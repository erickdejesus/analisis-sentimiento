2Pac	http://en.wikipedia.org/wiki/2pac
A. A. Milne	http://en.wikipedia.org/wiki/A._A._Milne
A. B. Guthrie	http://en.wikipedia.org/wiki/A._B._Guthrie
A. Bruce Bielaski	http://en.wikipedia.org/wiki/A._Bruce_Bielaski
A. E. Housman	http://en.wikipedia.org/wiki/A._E._Housman
A. E. van Vogt	http://en.wikipedia.org/wiki/A._E._van_Vogt
A. Edward Newton	http://en.wikipedia.org/wiki/A._Edward_Newton
A. J. Foyt	http://en.wikipedia.org/wiki/A._J._Foyt_IV
A. J. Liebling	http://en.wikipedia.org/wiki/A._J._Liebling
A. J. McLean	http://en.wikipedia.org/wiki/A._J._McLean
A. Jerrold Perenchio	http://en.wikipedia.org/wiki/A._Jerrold_Perenchio
A. L. Barker	http://en.wikipedia.org/wiki/A._L._Barker
A. Leon Higginbotham, Jr.	http://en.wikipedia.org/wiki/A._Leon_Higginbotham,_Jr.
A. N. Wilson	http://en.wikipedia.org/wiki/A._N._Wilson
A. Owsley Stanley	http://en.wikipedia.org/wiki/A._Owsley_Stanley
A. P. Giannini	http://en.wikipedia.org/wiki/A._P._Giannini
A. P. J. Kalam	http://en.wikipedia.org/wiki/A._P._J._Kalam
A. R. Ammons	http://en.wikipedia.org/wiki/A._R._Ammons
A. R. Radcliffe-Brown	http://en.wikipedia.org/wiki/A._R._Radcliffe-Brown
A. S. Byatt	http://en.wikipedia.org/wiki/A._S._Byatt
A. Whitney Brown	http://en.wikipedia.org/wiki/A._Whitney_Brown
A.D. Correll	http://en.wikipedia.org/wiki/A.D._%22Pete%22_Correll
Aage N. Bohr	http://en.wikipedia.org/wiki/Aage_N._Bohr
Aaliyah Dana Haughton	http://en.wikipedia.org/wiki/Aaliyah_Dana_Haughton
Aamir Khan	http://en.wikipedia.org/wiki/Aamir_Khan
Aaron Brown	http://en.wikipedia.org/wiki/Aaron_Brown
Aaron Burr	http://en.wikipedia.org/wiki/Aaron_Burr
Aaron Carter	http://en.wikipedia.org/wiki/Aaron_Carter
Aaron Cometbus	http://en.wikipedia.org/wiki/Aaron_Cometbus
Aaron Copland	http://en.wikipedia.org/wiki/Aaron_Copland
Aaron Eckhart	http://en.wikipedia.org/wiki/Aaron_Eckhart
Aaron Funk	http://en.wikipedia.org/wiki/Aaron_Funk
Aaron Hill	http://en.wikipedia.org/wiki/Aaron_Hill_(writer)
Aaron Klug	http://en.wikipedia.org/wiki/Aaron_Klug
Aaron Lewis	http://en.wikipedia.org/wiki/Aaron_Lewis
Aaron McGruder	http://en.wikipedia.org/wiki/Aaron_McGruder
Aaron Montgomery Ward	http://en.wikipedia.org/wiki/Aaron_Montgomery_Ward
Aaron Neville	http://en.wikipedia.org/wiki/Aaron_Neville
Aaron Schock	http://en.wikipedia.org/wiki/Aaron_Schock
Aaron Sorkin	http://en.wikipedia.org/wiki/Aaron_Sorkin
Aaron Spelling	http://en.wikipedia.org/wiki/Aaron_Spelling
Aaron Stanford	http://en.wikipedia.org/wiki/Aaron_Stanford
ABBA	http://en.wikipedia.org/wiki/Abba
Abba Eban	http://en.wikipedia.org/wiki/Abba_Eban
Abba Lerner	http://en.wikipedia.org/wiki/Abba_Lerner
Abbas El Fassi	http://en.wikipedia.org/wiki/Abbas_El_Fassi
Abbie Hoffman	http://en.wikipedia.org/wiki/Abbie_Hoffman
Abdel Aziz Rantisi	http://en.wikipedia.org/wiki/Abdel_Aziz_Rantisi
Abdelaziz Belkhadem	http://en.wikipedia.org/wiki/Abdelaziz_Belkhadem
Abdelaziz Bouteflika	http://en.wikipedia.org/wiki/Abdelaziz_Bouteflika
Abdelkader Taleb Oumar	http://en.wikipedia.org/wiki/Abdelkader_Taleb_Oumar
Abdou Soul� Elbak	http://en.wikipedia.org/wiki/Abdou_Soul%C3%A9_Elbak 
Abdoulaye Wade	http://en.wikipedia.org/wiki/Abdoulaye_Wade
Abdul Kalam	http://en.wikipedia.org/wiki/Abdul_Kalam
Abdul Qadeer Khan	http://en.wikipedia.org/wiki/Abdul_Qadeer_Khan
Abdul Qadir Bajamal	http://en.wikipedia.org/wiki/Abdul_Qadir_Bajamal
Abdul-Khalim Sadulayev	http://en.wikipedia.org/wiki/Abdul-Khalim_Sadulayev
Abdullah Ahmad Badawi	http://en.wikipedia.org/wiki/Abdullah_Ahmad_Badawi
Abdullah Azzam	http://en.wikipedia.org/wiki/Abdullah_Azzam
Abdullah G�l	http://en.wikipedia.org/wiki/Abdullah_G%C3%BCl
Abdullah ibn Khalifa Al Thani	http://en.wikipedia.org/wiki/Abdullah_ibn_Khalifa_Al_Thani
Abdullahi Yusuf	http://en.wikipedia.org/wiki/Abdullahi_Yusuf
Abdurrahman Wahid	http://en.wikipedia.org/wiki/Abdurrahman_Wahid
Abdus Salam	http://en.wikipedia.org/wiki/Abdus_Salam
Abe Fortas	http://en.wikipedia.org/wiki/Abe_Fortas
Abe Reles	http://en.wikipedia.org/wiki/Abe_Reles
Abe Vigoda	http://en.wikipedia.org/wiki/Abe_Vigoda
Abel Ferrara	http://en.wikipedia.org/wiki/Abel_Ferrara
Abel Gance	http://en.wikipedia.org/wiki/Abel_Gance
Abel Janszoon Tasman	http://en.wikipedia.org/wiki/Abel_Janszoon_Tasman
Abel Pacheco	http://en.wikipedia.org/wiki/Abel_Pacheco
Abhisit Vejjajiva	http://en.wikipedia.org/wiki/Abhisit_Vejjajiva
Abigail Adams	http://en.wikipedia.org/wiki/Abigail_Adams
Abigail Thernstrom	http://en.wikipedia.org/wiki/Abigail_Thernstrom
Abigail Van Buren	http://en.wikipedia.org/wiki/Abigail_Van_Buren
Abner Doubleday	http://en.wikipedia.org/wiki/Abner_Doubleday
Abner Haynes	http://en.wikipedia.org/wiki/Abner_Haynes
Abner Louima	http://en.wikipedia.org/wiki/Abner_Louima
Abolhassan Bani-Sadr	http://en.wikipedia.org/wiki/Abolhassan_Bani-Sadr
Abraham Benrubi	http://en.wikipedia.org/wiki/Abraham_Benrubi
Abraham de Moivre	http://en.wikipedia.org/wiki/Abraham_de_Moivre
Abraham Flexner	http://en.wikipedia.org/wiki/Abraham_Flexner
Abraham Gottlob Werner	http://en.wikipedia.org/wiki/Abraham_Gottlob_Werner
Abraham Lincoln	http://en.wikipedia.org/wiki/Abraham_Lincoln
Abraham Maslow	http://en.wikipedia.org/wiki/Abraham_Maslow
Abraham Ortelius	http://en.wikipedia.org/wiki/Abraham_Ortelius
Abraham Zapruder	http://en.wikipedia.org/wiki/Abraham_Zapruder
Abram Stevens Hewitt	http://en.wikipedia.org/wiki/Abram_Stevens_Hewitt
Abu Abbas	http://en.wikipedia.org/wiki/Abu_Abbas
Abu Bakar Bashir	http://en.wikipedia.org/wiki/Abu_Bakar_Bashir
Abu Faraj al-Libbi	http://en.wikipedia.org/wiki/Abu_Faraj_al-Libbi
Abu Hamza al-Masri	http://en.wikipedia.org/wiki/Abu_Hamza_al-Masri
Abu Mazen	http://en.wikipedia.org/wiki/Abu_Mazen
Abu Musab al-Zarqawi	http://en.wikipedia.org/wiki/Abu_Musab_al-Zarqawi
Abu Nidal	http://en.wikipedia.org/wiki/Abu_Nidal
Ace Frehley	http://en.wikipedia.org/wiki/Ace_Frehley
Ada Lovelace	http://en.wikipedia.org/wiki/Ada_Lovelace
Adalbert Stifter	http://en.wikipedia.org/wiki/Adalbert_Stifter
Adam Afriyie	http://en.wikipedia.org/wiki/Adam_Afriyie
Adam Ant	http://en.wikipedia.org/wiki/Adam_Ant
Adam Arkin	http://en.wikipedia.org/wiki/Adam_Arkin
Adam Baldwin	http://en.wikipedia.org/wiki/Adam_Baldwin
Adam Brody	http://en.wikipedia.org/wiki/Adam_Brody
Adam Carolla	http://en.wikipedia.org/wiki/Adam_Carolla
Adam Clayton	http://en.wikipedia.org/wiki/Adam_Clayton
Adam Clayton Powell	http://en.wikipedia.org/wiki/Adam_Clayton_Powell_IV_%28politician%29
Adam Clymer	http://en.wikipedia.org/wiki/Adam_Clymer
Adam Curry	http://en.wikipedia.org/wiki/Adam_Curry
Adam Duritz	http://en.wikipedia.org/wiki/Adam_Duritz
Adam Garcia	http://en.wikipedia.org/wiki/Adam_Garcia
Adam Gilchrist	http://en.wikipedia.org/wiki/Adam_Gilchrist
Adam Goldberg	http://en.wikipedia.org/wiki/Adam_Goldberg
Adam Holloway	http://en.wikipedia.org/wiki/Adam_Holloway
Adam Jones	http://en.wikipedia.org/wiki/Adam_Jones_%28musician%29
Adam Lamberg	http://en.wikipedia.org/wiki/Adam_Lamberg
Adam Levine	http://en.wikipedia.org/wiki/Adam_Levine
Adam Nagourney	http://en.wikipedia.org/wiki/Adam_Nagourney
Adam Osborne	http://en.wikipedia.org/wiki/Adam_Osborne
Adam Pascal	http://en.wikipedia.org/wiki/Adam_Pascal
Adam Posen	http://en.wikipedia.org/wiki/Adam_Posen
Adam Putnam	http://en.wikipedia.org/wiki/Adam_Putnam
Adam Rich	http://en.wikipedia.org/wiki/Adam_Rich
Adam Rickitt	http://en.wikipedia.org/wiki/Adam_Rickitt
Adam Sandler	http://en.wikipedia.org/wiki/Adam_Sandler
Adam Savage	http://en.wikipedia.org/wiki/Adam_Savage
Adam Schiff	http://en.wikipedia.org/wiki/Adam_Schiff
Adam Smith	http://en.wikipedia.org/wiki/Adam_Smith_%28politician%29
Adam Smith	http://en.wikipedia.org/wiki/Adam_Smith
Adam Weishaupt	http://en.wikipedia.org/wiki/Adam_Weishaupt
Adam West	http://en.wikipedia.org/wiki/Adam_West
Adele Addison	http://en.wikipedia.org/wiki/Adele_Addison
Adele Astaire	http://en.wikipedia.org/wiki/Adele_Astaire
Adele Mara	http://en.wikipedia.org/wiki/Adele_Mara
Adewale Akinnuoye-Agbaje	http://en.wikipedia.org/wiki/Adewale_Akinnuoye-Agbaje
Adil Abdul Mahdi	http://en.wikipedia.org/wiki/Adil_Abdul_Mahdi
Adlai E. Stevenson	http://en.wikipedia.org/wiki/Adlai_E._Stevenson_I
Adlai Stevenson	http://en.wikipedia.org/wiki/Adlai_Stevenson
Adnan Khashoggi	http://en.wikipedia.org/wiki/Adnan_Khashoggi
Adnan Pachachi	http://en.wikipedia.org/wiki/Adnan_Pachachi
Adnan Terzic	http://en.wikipedia.org/wiki/Adnan_Terzi%C4%87
Adolf Butenandt	http://en.wikipedia.org/wiki/Adolf_Butenandt
Adolf Eichmann	http://en.wikipedia.org/wiki/Adolf_Eichmann
Adolf Hitler	http://en.wikipedia.org/wiki/Adolf_Hitler
Adolf Loos	http://en.wikipedia.org/wiki/Adolf_Loos
Adolf von Baeyer	http://en.wikipedia.org/wiki/Adolf_von_Baeyer
Adolf Windaus	http://en.wikipedia.org/wiki/Adolf_Windaus
Adolfo Alix Jr.	http://en.wikipedia.org/wiki/Adolfo_Alix_Jr.
Adolfo Bioy Casares	http://en.wikipedia.org/wiki/Adolfo_Bioy_Casares
Adolfo Celi	http://en.wikipedia.org/wiki/Adolfo_Celi
Adolfo P�rez Esquivel	http://en.wikipedia.org/wiki/Adolfo_P%C3%A9rez_Esquivel
Adolph Dubs	http://en.wikipedia.org/wiki/Adolph_Dubs
Adolph Ochs	http://en.wikipedia.org/wiki/Adolph_Ochs
Adolphe Menjou	http://en.wikipedia.org/wiki/Adolphe_Menjou
Adolphe Muzito	http://en.wikipedia.org/wiki/Adolphe_Muzito
Adolphe Thiers	http://en.wikipedia.org/wiki/Adolphe_Thiers
Adolphe-William Bouguereau	http://en.wikipedia.org/wiki/Adolphe-William_Bouguereau
Adolphus Staton	http://en.wikipedia.org/wiki/Adolphus_Staton
Adoniram Judson	http://en.wikipedia.org/wiki/Adoniram_Judson
Adrian Adonis	http://en.wikipedia.org/wiki/Adrian_Adonis
Adrian Bailey	http://en.wikipedia.org/wiki/Adrian_Bailey
Adrian Belew	http://en.wikipedia.org/wiki/Adrian_Belew
Adrian Cronauer	http://en.wikipedia.org/wiki/Adrian_Cronauer
Adrian Edmondson	http://en.wikipedia.org/wiki/Adrian_Edmondson
Adrian Grenier	http://en.wikipedia.org/wiki/Adrian_Grenier
Adrian Lamo	http://en.wikipedia.org/wiki/Adrian_Lamo
Adrian Lyne	http://en.wikipedia.org/wiki/Adrian_Lyne
Adrian M. Smith	http://en.wikipedia.org/wiki/Adrian_M._Smith
Adrian Pasdar	http://en.wikipedia.org/wiki/Adrian_Pasdar
Adrian Paul	http://en.wikipedia.org/wiki/Adrian_Paul
Adrian Sanders	http://en.wikipedia.org/wiki/Adrian_Sanders
Adrian Zmed	http://en.wikipedia.org/wiki/Adrian_Zmed
Adriana Karembeu	http://en.wikipedia.org/wiki/Adriana_Karembeu
Adriana Lima	http://en.wikipedia.org/wiki/Adriana_Lima
Adrianne Curry	http://en.wikipedia.org/wiki/Adrianne_Curry
Adriano Castellesi	http://en.wikipedia.org/wiki/Adriano_Castellesi
Adrien Brody	http://en.wikipedia.org/wiki/Adrien_Brody
Adrien-Marie Legendre	http://en.wikipedia.org/wiki/Adrien-Marie_Legendre
Adrienne Albert	http://en.wikipedia.org/wiki/Adrienne_Albert
Adrienne Barbeau	http://en.wikipedia.org/wiki/Adrienne_Barbeau
Adrienne Rich	http://en.wikipedia.org/wiki/Adrienne_Rich
Aelius Aristides	http://en.wikipedia.org/wiki/Aelius_Aristides
Aelius Stilo	http://en.wikipedia.org/wiki/Aelius_Stilo
Aesop Rock	http://en.wikipedia.org/wiki/Aesop_Rock
Afrika Bambaataa	http://en.wikipedia.org/wiki/Afrika_Bambaataa
Agatha Christie	http://en.wikipedia.org/wiki/Agatha_Christie
Agim �eku	http://en.wikipedia.org/wiki/Agim_%C3%87eku
Agnes Bruckner	http://en.wikipedia.org/wiki/Agnes_Bruckner
Agnes de Mille	http://en.wikipedia.org/wiki/Agnes_de_Mille
Agnes Moorehead	http://en.wikipedia.org/wiki/Agnes_Moorehead
Agnes Strickland	http://en.wikipedia.org/wiki/Agnes_Strickland
Agnetha F�ltskog	http://en.wikipedia.org/wiki/Agnetha_F%C3%A4ltskog
Agostino Depretis	http://en.wikipedia.org/wiki/Agostino_Depretis
Agust�n de Iturbide	http://en.wikipedia.org/wiki/Agust%C3%ADn_de_Iturbide
Aharon Appelfeld	http://en.wikipedia.org/wiki/Aharon_Appelfeld
Ahmad Rashad	http://en.wikipedia.org/wiki/Ahmad_Rashad
Ahmad Tejan Kabbah	http://en.wikipedia.org/wiki/Ahmad_Tejan_Kabbah
Ahmed Abdallah Sambi	http://en.wikipedia.org/wiki/Ahmed_Abdallah_Sambi
Ahmed Ali	http://en.wikipedia.org/wiki/Ahmed_Ali
Ahmed Best	http://en.wikipedia.org/wiki/Ahmed_Best
Ahmed Chalabi	http://en.wikipedia.org/wiki/Ahmed_Chalabi
Ahmed H. Zewail	http://en.wikipedia.org/wiki/Ahmed_H._Zewail
Ahmed Khalfan Ghailani	http://en.wikipedia.org/wiki/Ahmed_Khalfan_Ghailani
Ahmed Nazif	http://en.wikipedia.org/wiki/Ahmed_Nazif
Ahmed Ouyahia	http://en.wikipedia.org/wiki/Ahmed_Ouyahia
Ahmed Qureia	http://en.wikipedia.org/wiki/Ahmed_Qurei
Ahmet Hadzipasic	http://en.wikipedia.org/wiki/Ahmet_Hadzipasic
Ahmet Necdet Sezer	http://en.wikipedia.org/wiki/Ahmet_Necdet_Sezer
Ahmet Zappa	http://en.wikipedia.org/wiki/Ahmet_Zappa
Aida Turturro	http://en.wikipedia.org/wiki/Aida_Turturro
Aidan Burley	http://en.wikipedia.org/wiki/Aidan_Burley
Aidan Quinn	http://en.wikipedia.org/wiki/Aidan_Quinn
Aigars Kalvitis	http://en.wikipedia.org/wiki/Aigars_Kalvitis
Aileen Quinn	http://en.wikipedia.org/wiki/Aileen_Quinn
Aileen Wuornos	http://en.wikipedia.org/wiki/Aileen_Wuornos
Aim� C�saire	http://en.wikipedia.org/wiki/Aim%C3%A9_C%C3%A9saire
Aimee Graham	http://en.wikipedia.org/wiki/Aimee_Graham
Aimee Mann	http://en.wikipedia.org/wiki/Aimee_Mann
Aimee Semple McPherson	http://en.wikipedia.org/wiki/Aimee_Semple_McPherson
Aires Ali	http://en.wikipedia.org/wiki/Aires_Ali
Aisha Tyler	http://en.wikipedia.org/wiki/Aisha_Tyler
Aishwarya Rai	http://en.wikipedia.org/wiki/Aishwarya_Rai
Ajay Devgan	http://en.wikipedia.org/wiki/Ajay_Devgan
Ajay Naidu	http://en.wikipedia.org/wiki/Ajay_Naidu
Akbar Abdi	http://en.wikipedia.org/wiki/Akbar_Abdi
Akbar Hashemi Rafsanjani	http://en.wikipedia.org/wiki/Akbar_Hashemi_Rafsanjani
Akbar the Great	http://en.wikipedia.org/wiki/Akbar_the_Great
Akhmad Kadyrov	http://en.wikipedia.org/wiki/Akhmad_Kadyrov
Aki Aleong	http://en.wikipedia.org/wiki/Aki_Aleong
Akil Akilov	http://en.wikipedia.org/wiki/Akil_Akilov
Akio Morita	http://en.wikipedia.org/wiki/Akio_Morita
Akira Kurosawa	http://en.wikipedia.org/wiki/Akira_Kurosawa
Akshay Kumar	http://en.wikipedia.org/wiki/Akshay_Kumar
Akshaye Khanna	http://en.wikipedia.org/wiki/Akshaye_Khanna
Al Capone	http://en.wikipedia.org/wiki/Al_Capone
Al Capp	http://en.wikipedia.org/wiki/Al_Capp
Al D'Amato	http://en.wikipedia.org/wiki/Al_D%27Amato
Al Davis	http://en.wikipedia.org/wiki/Al_Davis
Al Di Meola	http://en.wikipedia.org/wiki/Al_Di_Meola
Al Franken	http://en.wikipedia.org/wiki/Al_Franken
Al Goldstein	http://en.wikipedia.org/wiki/Al_Goldstein
Al Gore	http://en.wikipedia.org/wiki/Al_Gore
Al Green	http://en.wikipedia.org/wiki/Al_Green_%28Texas%29
Al Green	http://en.wikipedia.org/wiki/Al_Green
Al Hirschfeld	http://en.wikipedia.org/wiki/Al_Hirschfeld
Al Hirt	http://en.wikipedia.org/wiki/Al_Hirt
Al Hunt	http://en.wikipedia.org/wiki/Al_Hunt
Al Jarreau	http://en.wikipedia.org/wiki/Al_Jarreau
Al Jolson	http://en.wikipedia.org/wiki/Al_Jolson
Al Jourgensen	http://en.wikipedia.org/wiki/Al_Jourgensen
Al Kaline	http://en.wikipedia.org/wiki/Al_Kaline
Al Lewis	http://en.wikipedia.org/wiki/Al_Lewis_%28actor%29
Al Lopez	http://en.wikipedia.org/wiki/Al_Lopez
Al McCandless	http://en.wikipedia.org/wiki/Al_McCandless
Al Michaels	http://en.wikipedia.org/wiki/Al_Michaels
Al Molinaro	http://en.wikipedia.org/wiki/Al_Molinaro
Al Pacino	http://en.wikipedia.org/wiki/Al_Pacino
Al Reynolds	http://en.wikipedia.org/wiki/Al_Reynolds
Al Roker	http://en.wikipedia.org/wiki/Al_Roker
Al Sapienza	http://en.wikipedia.org/wiki/Al_Sapienza
Al Sharpton	http://en.wikipedia.org/wiki/Al_Sharpton
Al Simmons	http://en.wikipedia.org/wiki/Al_Simmons
Al Stewart	http://en.wikipedia.org/wiki/Al_Stewart
Al Swift	http://en.wikipedia.org/wiki/Al_Swift
Al Unser, Jr.	http://en.wikipedia.org/wiki/Al_Unser,_Jr.
Al Unser, Sr.	http://en.wikipedia.org/wiki/Al_Unser,_Sr.
Alain Chartier	http://en.wikipedia.org/wiki/Alain_Chartier
Alain Delon	http://en.wikipedia.org/wiki/Alain_Delon
Alain J. P. Belda	http://en.wikipedia.org/wiki/Alain_J._P._Belda
Alain Jupp�	http://en.wikipedia.org/wiki/Alain_Jupp%C3%A9
Alain Locke	http://en.wikipedia.org/wiki/Alain_Locke
Alain Ren� Lesage	http://en.wikipedia.org/wiki/Alain_Ren%C3%A9_Lesage
Alain Robbe-Grillet	http://en.wikipedia.org/wiki/Alain_Robbe-Grillet
Alain Robert	http://en.wikipedia.org/wiki/Alain_Robert
Alan Alda	http://en.wikipedia.org/wiki/Alan_Alda
Alan Arkin	http://en.wikipedia.org/wiki/Alan_Arkin
Alan Autry	http://en.wikipedia.org/wiki/Alan_Autry
Alan B. Mollohan	http://en.wikipedia.org/wiki/Alan_B._Mollohan
Alan Ball	http://en.wikipedia.org/wiki/Alan_Ball_%28screenwriter%29
Alan Ball	http://en.wikipedia.org/wiki/Allan_Ball
Alan Bates	http://en.wikipedia.org/wiki/Alan_Bates
Alan Bean	http://en.wikipedia.org/wiki/Alan_Bean
Alan Beith	http://en.wikipedia.org/wiki/Alan_Beith
Alan Bennett	http://en.wikipedia.org/wiki/Alan_Bennett
Alan Bullock	http://en.wikipedia.org/wiki/Alan_Bullock
Alan Campbell	http://en.wikipedia.org/wiki/Alan_Campbell_%28writer%29
Alan Colmes	http://en.wikipedia.org/wiki/Alan_Colmes
Alan Cox	http://en.wikipedia.org/wiki/Alan_Cox
Alan Cranston	http://en.wikipedia.org/wiki/Alan_Cranston
Alan Cumming	http://en.wikipedia.org/wiki/Alan_Cumming
Alan Dale	http://en.wikipedia.org/wiki/Alan_Dale
Alan Dean Foster	http://en.wikipedia.org/wiki/Alan_Dean_Foster
Alan Dershowitz	http://en.wikipedia.org/wiki/Alan_Dershowitz
Alan Dugan	http://en.wikipedia.org/wiki/Alan_Dugan
Alan Duncan	http://en.wikipedia.org/wiki/Alan_Duncan
Alan Freed	http://en.wikipedia.org/wiki/Alan_Freed
Alan G. MacDiarmid	http://en.wikipedia.org/wiki/Alan_G._MacDiarmid
Alan Garc�a	http://en.wikipedia.org/wiki/Alan_Garc%C3%ADa
Alan Gowen	http://en.wikipedia.org/wiki/Alan_Gowen
Alan Grayson	http://en.wikipedia.org/wiki/Alan_Grayson
Alan Greenspan	http://en.wikipedia.org/wiki/Alan_Greenspan
Alan Hale, Jr.	http://en.wikipedia.org/wiki/Alan_Hale,_Jr.
Alan Hale, Sr.	http://en.wikipedia.org/wiki/Alan_Hale,_Sr.
Alan Hansen	http://en.wikipedia.org/wiki/Alan_Hansen
Alan Haselhurst	http://en.wikipedia.org/wiki/Alan_Haselhurst
Alan J. Dixon	http://en.wikipedia.org/wiki/Alan_J._Dixon
Alan J. Heeger	http://en.wikipedia.org/wiki/Alan_J._Heeger
Alan J. Lacy	http://en.wikipedia.org/wiki/Alan_J._Lacy
Alan J. Pakula	http://en.wikipedia.org/wiki/Alan_J._Pakula
Alan Jackson	http://en.wikipedia.org/wiki/Alan_Jackson
Alan Johnson	http://en.wikipedia.org/wiki/Alan_Johnson
Alan K. Simpson	http://en.wikipedia.org/wiki/Alan_K._Simpson
Alan Kay	http://en.wikipedia.org/wiki/Alan_Kay
Alan Keen	http://en.wikipedia.org/wiki/Alan_Keen
Alan Keyes	http://en.wikipedia.org/wiki/Alan_Keyes
Alan King	http://en.wikipedia.org/wiki/Alan_King_%28comedian%29
Alan L. Boeckmann	http://en.wikipedia.org/wiki/Alan_L._Boeckmann
Alan Ladd	http://en.wikipedia.org/wiki/Alan_Ladd
Alan Lomax	http://en.wikipedia.org/wiki/Alan_Lomax
Alan Meale	http://en.wikipedia.org/wiki/Alan_Meale
Alan Miller	http://en.wikipedia.org/wiki/Alan_Miller_%28game_designer%29
Alan Minter	http://en.wikipedia.org/wiki/Alan_Minter
Alan Mollohan	http://en.wikipedia.org/wiki/Alan_Mollohan
Alan Moore	http://en.wikipedia.org/wiki/Alan_Moore
Alan Moulder	http://en.wikipedia.org/wiki/Alan_Moulder
Alan Mowbray	http://en.wikipedia.org/wiki/Alan_Mowbray
Alan Myerson	http://en.wikipedia.org/wiki/Alan_Myerson
Alan Napier	http://en.wikipedia.org/wiki/Alan_Napier
Alan Osmond	http://en.wikipedia.org/wiki/Alan_Osmond
Alan Page	http://en.wikipedia.org/wiki/Alan_Page
Alan Parker	http://en.wikipedia.org/wiki/Alan_Parker
Alan Parsons	http://en.wikipedia.org/wiki/Alan_Parsons
Alan Paton	http://en.wikipedia.org/wiki/Alan_Paton
Alan Reed	http://en.wikipedia.org/wiki/Alan_Reed
Alan Reid	http://en.wikipedia.org/wiki/Alan_Reed
Alan Rickman	http://en.wikipedia.org/wiki/Alan_Rickman
Alan Ruck	http://en.wikipedia.org/wiki/Alan_Ruck
Alan Rudolph	http://en.wikipedia.org/wiki/Alan_Rudolph
Alan S. Boyd	http://en.wikipedia.org/wiki/Alan_S._Boyd
Alan Shearer	http://en.wikipedia.org/wiki/Alan_Shearer
Alan Shepard	http://en.wikipedia.org/wiki/Alan_Shepard
Alan Shugart	http://en.wikipedia.org/wiki/Alan_Shugart
Alan Sillitoe	http://en.wikipedia.org/wiki/Alan_Sillitoe
Alan Simpson	http://en.wikipedia.org/wiki/Alan_Simpson_%28politician%29
Alan Sokal	http://en.wikipedia.org/wiki/Alan_Sokal
Alan Thicke	http://en.wikipedia.org/wiki/Alan_Thicke
Alan Turing	http://en.wikipedia.org/wiki/Alan_Turing
Alan Vega	http://en.wikipedia.org/wiki/Alan_Vega
Alan Watson Steelman	http://en.wikipedia.org/wiki/Alan_Watson
Alan Wheat	http://en.wikipedia.org/wiki/Alan_Wheat
Alan White	http://en.wikipedia.org/wiki/Alan_White_%28Yes_drummer%29
Alan Whitehead	http://en.wikipedia.org/wiki/Alan_Whitehead
Alan Young	http://en.wikipedia.org/wiki/Alan_Young
Alanis Morissette	http://en.wikipedia.org/wiki/Alanis_Morissette
Alannah Myles	http://en.wikipedia.org/wiki/Alannah_Myles
Alaric I	http://en.wikipedia.org/wiki/Alaric_I
Alasdair McDonnell	http://en.wikipedia.org/wiki/Alasdair_McDonnell
Alastair Sim	http://en.wikipedia.org/wiki/Alastair_Sim
Alban Berg	http://en.wikipedia.org/wiki/Alban_Berg
Alban Butler	http://en.wikipedia.org/wiki/Alban_Butler
Alben W. Barkley	http://en.wikipedia.org/wiki/Alben_W._Barkley
Alberico Gentili	http://en.wikipedia.org/wiki/Alberico_Gentili
Albert A. Michelson	http://en.wikipedia.org/wiki/Albert_A._Michelson
Albert Anastasia	http://en.wikipedia.org/wiki/Albert_Anastasia
Albert Ayler	http://en.wikipedia.org/wiki/Albert_Ayler
Albert Bassermann	http://en.wikipedia.org/wiki/Albert_Bassermann
Albert Brooks	http://en.wikipedia.org/wiki/Albert_Brooks
Albert Camille Vital	http://en.wikipedia.org/wiki/Albert_Camille_Vital
Albert Camus	http://en.wikipedia.org/wiki/Albert_Camus
Albert Dekker	http://en.wikipedia.org/wiki/Albert_Dekker
Albert Einstein	http://en.wikipedia.org/wiki/Albert_Einstein
Albert Finney	http://en.wikipedia.org/wiki/Albert_Finney
Albert Fish	http://en.wikipedia.org/wiki/Albert_Fish
Albert G. Bustamante	http://en.wikipedia.org/wiki/Albert_G._Bustamante
Albert Gallatin	http://en.wikipedia.org/wiki/Albert_Gallatin
Albert Gobat	http://en.wikipedia.org/wiki/Albert_Gobat
Albert Goldbarth	http://en.wikipedia.org/wiki/Albert_Goldbarth
Albert Hofmann	http://en.wikipedia.org/wiki/Albert_Hofmann
Albert Hughes	http://en.wikipedia.org/wiki/Albert_Hughes
Albert I	http://en.wikipedia.org/wiki/Albert_I_of_Belgium
Albert II	http://en.wikipedia.org/wiki/Albert_II_of_Belgium
Albert Jay Nock	http://en.wikipedia.org/wiki/Albert_Jay_Nock
Albert King	http://en.wikipedia.org/wiki/Albert_King
Albert L. Murray	http://en.wikipedia.org/wiki/Albert_L._Murray
Albert Lutuli	http://en.wikipedia.org/wiki/Albert_Lutuli
Albert Maltz	http://en.wikipedia.org/wiki/Albert_Maltz
Albert Maysles	http://en.wikipedia.org/wiki/Albert_Maysles
Albert Moore	http://en.wikipedia.org/wiki/Albert_Joseph_Moore
Albert Owen	http://en.wikipedia.org/wiki/Albert_Owen
Albert Pinkham Ryder	http://en.wikipedia.org/wiki/Albert_Pinkham_Ryder
Albert Pintat	http://en.wikipedia.org/wiki/Albert_Pintat
Albert Pujols	http://en.wikipedia.org/wiki/Albert_Pujols
Albert Pyun	http://en.wikipedia.org/wiki/Albert_Pyun
Albert R. Broccoli	http://en.wikipedia.org/wiki/Albert_R._Broccoli
Albert Reynolds	http://en.wikipedia.org/wiki/Albert_Reynolds
Albert Sabin	http://en.wikipedia.org/wiki/Albert_Sabin
Albert Schweitzer	http://en.wikipedia.org/wiki/Albert_Schweitzer
Albert Sidney Johnston	http://en.wikipedia.org/wiki/Albert_Sidney_Johnston
Albert Speer	http://en.wikipedia.org/wiki/Albert_Speer
Albert V. Casey	http://en.wikipedia.org/wiki/Albert_Vincent_Casey
Albert Wallace Hull	http://en.wikipedia.org/wiki/Albert_Wallace_Hull
Albert Wohlstetter	http://en.wikipedia.org/wiki/Albert_Wohlstetter
Albert Wynn	http://en.wikipedia.org/wiki/Albert_Wynn
Alberta Hunter	http://en.wikipedia.org/wiki/Alberta_Hunter
Alberto Acosta	http://en.wikipedia.org/wiki/Alberto_Acosta
Alberto Fujimori	http://en.wikipedia.org/wiki/Alberto_Fujimori
Alberto Giacometti	http://en.wikipedia.org/wiki/Alberto_Giacometti
Alberto Gonzales	http://en.wikipedia.org/wiki/Alberto_Gonzales
Alberto Moravia	http://en.wikipedia.org/wiki/Alberto_Moravia
Alberto Vargas	http://en.wikipedia.org/wiki/Alberto_Vargas
Albio Sires	http://en.wikipedia.org/wiki/Albio_Sires
Albrecht Altdorfer	http://en.wikipedia.org/wiki/Albrecht_Altdorfer
Albrecht D�rer	http://en.wikipedia.org/wiki/Albrecht_D%C3%BCrer
Albrecht von Haller	http://en.wikipedia.org/wiki/Albrecht_von_Haller
Albrecht von Wallenstein	http://en.wikipedia.org/wiki/Albrecht_von_Wallenstein
Alcee Hastings	http://en.wikipedia.org/wiki/Alcee_Hastings
Aldo Leopold	http://en.wikipedia.org/wiki/Aldo_Leopold
Aldo Moro	http://en.wikipedia.org/wiki/Aldo_Moro
Aldo Ray	http://en.wikipedia.org/wiki/Aldo_Ray
Aldous Huxley	http://en.wikipedia.org/wiki/Aldous_Huxley
Aldrich Ames	http://en.wikipedia.org/wiki/Aldrich_Ames
Aldus Manutius	http://en.wikipedia.org/wiki/Aldus_Manutius
Alec Baldwin	http://en.wikipedia.org/wiki/Alec_Baldwin
Alec Douglas-Home	http://en.wikipedia.org/wiki/Alec_Douglas-Home
Alec Empire	http://en.wikipedia.org/wiki/Alec_Empire
Alec Guinness	http://en.wikipedia.org/wiki/Alec_Guinness
Alec Shelbrooke	http://en.wikipedia.org/wiki/Alec_Shelbrooke
Alec Waugh	http://en.wikipedia.org/wiki/Alec_Waugh
Aleister Crowley	http://en.wikipedia.org/wiki/Aleister_Crowley
Alejandro Sanz	http://en.wikipedia.org/wiki/Alejandro_Sanz
Alejandro Toledo	http://en.wikipedia.org/wiki/Alejandro_Toledo
Aleksander Bovin	http://en.wikipedia.org/wiki/Alexander_Bovin
Aleksander Kwasniewski	http://en.wikipedia.org/wiki/Aleksander_Kwasniewski
Aleksandr Borodin	http://en.wikipedia.org/wiki/Aleksandr_Borodin
Aleksandr Glazunov	http://en.wikipedia.org/wiki/Aleksandr_Glazunov
Aleksandr Lukashenko	http://en.wikipedia.org/wiki/Aleksandr_Lukashenko
Aleksandr M. Prokhorov	http://en.wikipedia.org/wiki/Aleksandr_M._Prokhorov
Aleksandr Pushkin	http://en.wikipedia.org/wiki/Aleksandr_Pushkin
Aleksandr Scriabin	http://en.wikipedia.org/wiki/Aleksandr_Scriabin
Aleksandr Sumarokov	http://en.wikipedia.org/wiki/Aleksandr_Sumarokov
Alessandro Farnese	http://en.wikipedia.org/wiki/Alessandro_Farnese,_Duke_of_Parma_and_Piacenza
Alessandro Manzoni	http://en.wikipedia.org/wiki/Alessandro_Manzoni
Alessandro Scarlatti	http://en.wikipedia.org/wiki/Alessandro_Scarlatti
Alessandro Stradella	http://en.wikipedia.org/wiki/Alessandro_Stradella
Alessandro Tassoni	http://en.wikipedia.org/wiki/Alessandro_Tassoni
Alessandro Volta	http://en.wikipedia.org/wiki/Alessandro_Volta
Alesso Baldovinetti	http://en.wikipedia.org/wiki/Alesso_Baldovinetti
Alex Barris	http://en.wikipedia.org/wiki/Alex_Barris
Alex Borstein	http://en.wikipedia.org/wiki/Alex_Borstein
Alex Chilton	http://en.wikipedia.org/wiki/Alex_Chilton
Alex Cord	http://en.wikipedia.org/wiki/Alex_Cord
Alex Cunningham	http://en.wikipedia.org/wiki/Alex_Cunningham
Alex Haley	http://en.wikipedia.org/wiki/Alex_Haley
Alex James	http://en.wikipedia.org/wiki/Alex_James_%28musician%29
Alex Jones	http://en.wikipedia.org/wiki/Alex_Jones_%28radio_host%29
Alex Kapranos	http://en.wikipedia.org/wiki/Alex_Kapranos
Alex Karras	http://en.wikipedia.org/wiki/Alex_Karras
Alex Kingston	http://en.wikipedia.org/wiki/Alex_Kingston
Alex Lifeson	http://en.wikipedia.org/wiki/Alex_Lifeson
Alex McMillan	http://en.wikipedia.org/wiki/Alex_McMillan
Alex Patterson	http://en.wikipedia.org/wiki/Alex_Patterson
Alex Penelas	http://en.wikipedia.org/wiki/Alex_Penelas
Alex Rocco	http://en.wikipedia.org/wiki/Alex_Rocco
Alex Rodriguez	http://en.wikipedia.org/wiki/Alex_Rodriguez
Alex Toth	http://en.wikipedia.org/wiki/Alex_Toth
Alex Trebek	http://en.wikipedia.org/wiki/Alex_Trebek
Alex Van Halen	http://en.wikipedia.org/wiki/Alex_Van_Halen
Alex Winter	http://en.wikipedia.org/wiki/Alex_Winter
Alexa Vega	http://en.wikipedia.org/wiki/Alexa_Vega
Alexander A. Vandegrift	http://en.wikipedia.org/wiki/Alexander_A._Vandegrift
Alexander Ankvab	http://en.wikipedia.org/wiki/Alexander_Ankvab
Alexander Bain	http://en.wikipedia.org/wiki/Alexander_Bain
Alexander Bickel	http://en.wikipedia.org/wiki/Alexander_Bickel
Alexander Blok	http://en.wikipedia.org/wiki/Alexander_Blok
Alexander Calder	http://en.wikipedia.org/wiki/Alexander_Calder
Alexander Cockburn	http://en.wikipedia.org/wiki/Alexander_Cockburn
Alexander Cruden	http://en.wikipedia.org/wiki/Alexander_Cruden
Alexander Downer	http://en.wikipedia.org/wiki/Alexander_Downer
Alexander Dubcek	http://en.wikipedia.org/wiki/Alexander_Dubcek
Alexander Fleming	http://en.wikipedia.org/wiki/Alexander_Fleming
Alexander Godunov	http://en.wikipedia.org/wiki/Alexander_Godunov
Alexander Gordon Laing	http://en.wikipedia.org/wiki/Alexander_Gordon_Laing
Alexander Graham Bell	http://en.wikipedia.org/wiki/Alexander_Graham_Bell
Alexander Haig	http://en.wikipedia.org/wiki/Alexander_Haig
Alexander Hamilton	http://en.wikipedia.org/wiki/Alexander_Hamilton
Alexander Hamilton Stephens	http://en.wikipedia.org/wiki/Alexander_Hamilton_Stephens
Alexander Kerensky	http://en.wikipedia.org/wiki/Alexander_Kerensky
Alexander Korda	http://en.wikipedia.org/wiki/Alexander_Korda
Alexander Lukashenko	http://en.wikipedia.org/wiki/Alexander_Lukashenko
Alexander Luria	http://en.wikipedia.org/wiki/Alexander_Luria
Alexander M. Poniatoff	http://en.wikipedia.org/wiki/Alexander_M._Poniatoff
Alexander Mackendrick	http://en.wikipedia.org/wiki/Alexander_Mackendrick
Alexander Mackenzie	http://en.wikipedia.org/wiki/Alexander_Mackenzie
Alexander Payne	http://en.wikipedia.org/wiki/Alexander_Payne
Alexander Pope	http://en.wikipedia.org/wiki/Alexander_Pope
Alexander R. Todd	http://en.wikipedia.org/wiki/Alexander_R._Todd
Alexander Siddig	http://en.wikipedia.org/wiki/Alexander_Siddig
Alexander Solzhenitsyn	http://en.wikipedia.org/wiki/Alexander_Solzhenitsyn
Alexander Suvorov	http://en.wikipedia.org/wiki/Alexander_Suvorov
Alexander the Great	http://en.wikipedia.org/wiki/Alexander_the_Great
Alexander Trowbridge	http://en.wikipedia.org/wiki/Alexander_Trowbridge
Alexander von Schlippenbach	http://en.wikipedia.org/wiki/Alexander_von_Schlippenbach
Alexander Woollcott	http://en.wikipedia.org/wiki/Alexander_Woollcott
Alexandra Hedison	http://en.wikipedia.org/wiki/Alexandra_Hedison
Alexandra Paul	http://en.wikipedia.org/wiki/Alexandra_Paul
Alexandra Ripley	http://en.wikipedia.org/wiki/Alexandra_Ripley
Alexandre Decamps	http://en.wikipedia.org/wiki/Alexandre_Decamps
Alexandre Dumas fils	http://en.wikipedia.org/wiki/Alexandre_Dumas_fils
Alexandre Dumas p�re	http://en.wikipedia.org/wiki/Alexandre_Dumas_p%C3%A8re
Alexei A. Abrikosov	http://en.wikipedia.org/wiki/Alexei_Alexeyevich_Abrikosov
Alexei Kosygin	http://en.wikipedia.org/wiki/Alexei_Kosygin
Alexei Leonov	http://en.wikipedia.org/wiki/Alexei_Leonov
Alexey Pajitnov	http://en.wikipedia.org/wiki/Alexey_Pajitnov
Alexi Laiho	http://en.wikipedia.org/wiki/Alexi_Laiho
Alexis Arquette	http://en.wikipedia.org/wiki/Alexis_Arquette
Alexis Bledel	http://en.wikipedia.org/wiki/Alexis_Bledel
Alexis de Tocqueville	http://en.wikipedia.org/wiki/Alexis_de_Tocqueville
Alexis Denisof	http://en.wikipedia.org/wiki/Alexis_Denisof
Alexis Herman	http://en.wikipedia.org/wiki/Alexis_Herman
Alexis Korner	http://en.wikipedia.org/wiki/Alexis_Korner
Alexis Smith	http://en.wikipedia.org/wiki/Alexis_Smith
Alf Landon	http://en.wikipedia.org/wiki/Alf_Landon
Alferd Packer	http://en.wikipedia.org/wiki/Alferd_Packer
Alfonse M. D'Amato	http://en.wikipedia.org/wiki/Alfonse_M._D%27Amato
Alfonso Garc�a Robles	http://en.wikipedia.org/wiki/Alfonso_Garc%C3%ADa_Robles
Alfonso Ribeiro	http://en.wikipedia.org/wiki/Alfonso_Ribeiro
Alfre Woodard	http://en.wikipedia.org/wiki/Alfre_Woodard
Alfred A. Knopf	http://en.wikipedia.org/wiki/Alfred_A._Knopf,_Sr.
Alfred Adler	http://en.wikipedia.org/wiki/Alfred_Adler
Alfred Austin	http://en.wikipedia.org/wiki/Alfred_Austin
Alfred Bester	http://en.wikipedia.org/wiki/Alfred_Bester
Alfred Chandler	http://en.wikipedia.org/wiki/Alfred_D._Chandler,_Jr.
Alfred Chester	http://en.wikipedia.org/wiki/Alfred_Chester
Alfred Cornu	http://en.wikipedia.org/wiki/Alfred_Cornu
Alfred de Musset	http://en.wikipedia.org/wiki/Alfred_de_Musset
Alfred de Vigny	http://en.wikipedia.org/wiki/Alfred_de_Vigny
Alfred Dreyfus	http://en.wikipedia.org/wiki/Alfred_Dreyfus
Alfred E. Smith	http://en.wikipedia.org/wiki/Alfred_E._Smith
Alfred Eisenstaedt	http://en.wikipedia.org/wiki/Alfred_Eisenstaedt
Alfred Fried	http://en.wikipedia.org/wiki/Alfred_Fried
Alfred Hitchcock	http://en.wikipedia.org/wiki/Alfred_Hitchcock
Alfred Jarry	http://en.wikipedia.org/wiki/Alfred_Jarry
Alfred Jodl	http://en.wikipedia.org/wiki/Alfred_Jodl
Alfred Kastler	http://en.wikipedia.org/wiki/Alfred_Kastler
Alfred Kazin	http://en.wikipedia.org/wiki/Alfred_Kazin
Alfred Kinsey	http://en.wikipedia.org/wiki/Alfred_Kinsey
Alfred Kreymborg	http://en.wikipedia.org/wiki/Alfred_Kreymborg
Alfred Kroeber	http://en.wikipedia.org/wiki/Alfred_Kroeber
Alfred Lord Tennyson	http://en.wikipedia.org/wiki/Alfred_Lord_Tennyson
Alfred Lunt	http://en.wikipedia.org/wiki/Alfred_Lunt
Alfred Moisiu	http://en.wikipedia.org/wiki/Alfred_Moisiu
Alfred Molina	http://en.wikipedia.org/wiki/Alfred_Molina
Alfred Newman	http://en.wikipedia.org/wiki/Alfred_Newman
Alfred Nobel	http://en.wikipedia.org/wiki/Alfred_Nobel
Alfred North Whitehead	http://en.wikipedia.org/wiki/Alfred_North_Whitehead
Alfred P. Murrah	http://en.wikipedia.org/wiki/Alfred_P._Murrah
Alfred P. Sloan	http://en.wikipedia.org/wiki/Alfred_P._Sloan
Alfred P. Swineford	http://en.wikipedia.org/wiki/Alfred_P._Swineford
Alfred Peet	http://en.wikipedia.org/wiki/Alfred_Peet
Alfred R. Berkeley III	http://en.wikipedia.org/wiki/Alfred_Berkeley
Alfred Rosenberg	http://en.wikipedia.org/wiki/Alfred_Rosenberg
Alfred Russel Wallace	http://en.wikipedia.org/wiki/Alfred_Russel_Wallace
Alfred Stevens	http://en.wikipedia.org/wiki/Alfred_Stevens_%28sculptor%29
Alfred Stieglitz	http://en.wikipedia.org/wiki/Alfred_Stieglitz
Alfred Tarski	http://en.wikipedia.org/wiki/Alfred_Tarski
Alfred von Tirpitz	http://en.wikipedia.org/wiki/Alfred_von_Tirpitz
Alfred Werner	http://en.wikipedia.org/wiki/Alfred_Werner
Alfredo Casella	http://en.wikipedia.org/wiki/Alfredo_Casella
Alfredo Di Stefano	http://en.wikipedia.org/wiki/Alfredo_Di_Stefano
Alfredo Palacio	http://en.wikipedia.org/wiki/Alfredo_Palacio
Alfredo Stroessner	http://en.wikipedia.org/wiki/Alfredo_Stroessner
Alfried Krupp	http://en.wikipedia.org/wiki/Alfried_Krupp
Alger Hiss	http://en.wikipedia.org/wiki/Alger_Hiss
Algernon Charles Swinburne	http://en.wikipedia.org/wiki/Algernon_Charles_Swinburne
Algernon Sidney	http://en.wikipedia.org/wiki/Algernon_Sidney
Algirdas Brazauskas	http://en.wikipedia.org/wiki/Algirdas_Brazauskas
Ali Abassi	http://en.wikipedia.org/wiki/Ali_Abassi
Ali Abdullah Saleh	http://en.wikipedia.org/wiki/Ali_Abdullah_Saleh
Ali Bongo Ondimba	http://en.wikipedia.org/wiki/Ali_Bongo_Ondimba
Ali Farka Tour�	http://en.wikipedia.org/wiki/Ali_Farka_Tour%C3%A9
Ali G	http://en.wikipedia.org/wiki/Ali_G
Ali Khamenei	http://en.wikipedia.org/wiki/Ali_Khamenei
Ali Landry	http://en.wikipedia.org/wiki/Ali_Landry
Ali Larter	http://en.wikipedia.org/wiki/Ali_Larter
Ali MacGraw	http://en.wikipedia.org/wiki/Ali_MacGraw
Ali Muhammad Ghedi	http://en.wikipedia.org/wiki/Ali_Muhammad_Ghedi
Ali Muhammad Mujawar	http://en.wikipedia.org/wiki/Ali_Muhammad_Mujawar
Alia Shawkat	http://en.wikipedia.org/wiki/Alia_Shawkat
Alice B. Toklas	http://en.wikipedia.org/wiki/Alice_B._Toklas
Alice Brady	http://en.wikipedia.org/wiki/Alice_Brady
Alice Cooper	http://en.wikipedia.org/wiki/Alice_Cooper
Alice Dunbar-Nelson	http://en.wikipedia.org/wiki/Alice_Dunbar-Nelson
Alice Faye	http://en.wikipedia.org/wiki/Alice_Faye
Alice Grant Rosman	http://en.wikipedia.org/wiki/Alice_Grant_Rosman
Alice Guy	http://en.wikipedia.org/wiki/Alice_Guy
Alice Hegan Rice	http://en.wikipedia.org/wiki/Alice_Hegan_Rice
Alice Hoffman	http://en.wikipedia.org/wiki/Alice_Hoffman
Alice Munro	http://en.wikipedia.org/wiki/Alice_Munro
Alice Paul	http://en.wikipedia.org/wiki/Alice_Paul
Alice Rivlin	http://en.wikipedia.org/wiki/Alice_Rivlin
Alice Roosevelt Longworth	http://en.wikipedia.org/wiki/Alice_Roosevelt_Longworth
Alice Walker	http://en.wikipedia.org/wiki/Alice_Walker
Alice Walton	http://en.wikipedia.org/wiki/Alice_Walton
Alicia Goranson	http://en.wikipedia.org/wiki/Alicia_Goranson
Alicia Keys	http://en.wikipedia.org/wiki/Alicia_Keys
Alicia Silverstone	http://en.wikipedia.org/wiki/Alicia_Silverstone
Alicia Witt	http://en.wikipedia.org/wiki/Alicia_Witt
Alida Valli	http://en.wikipedia.org/wiki/Alida_Valli
Alison Arngrim	http://en.wikipedia.org/wiki/Alison_Arngrim
Alison Bechdel	http://en.wikipedia.org/wiki/Alison_Bechdel
Alison Eastwood	http://en.wikipedia.org/wiki/Alison_Eastwood
Alison Krauss	http://en.wikipedia.org/wiki/Alison_Krauss
Alison Lohman	http://en.wikipedia.org/wiki/Alison_Lohman
Alison Lurie	http://en.wikipedia.org/wiki/Alison_Lurie
Alison McGovern	http://en.wikipedia.org/wiki/Alison_McGovern
Alison Moyet	http://en.wikipedia.org/wiki/Alison_Moyet
Alison Seabeck	http://en.wikipedia.org/wiki/Alison_Seabeck
Alistair Burt	http://en.wikipedia.org/wiki/Alistair_Burt
Alistair Carmichael	http://en.wikipedia.org/wiki/Alistair_Carmichael
Alistair Cooke	http://en.wikipedia.org/wiki/Alistair_Cooke
Alistair Darling	http://en.wikipedia.org/wiki/Alistair_Darling
Allan Ahlberg	http://en.wikipedia.org/wiki/Allan_Ahlberg
Allan Albert	http://en.wikipedia.org/wiki/Allan_Albert
Allan Arbus	http://en.wikipedia.org/wiki/Allan_Arbus
Allan Bloom	http://en.wikipedia.org/wiki/Allan_Bloom
Allan Dwan	http://en.wikipedia.org/wiki/Allan_Dwan
Allan Gurganus	http://en.wikipedia.org/wiki/Allan_Gurganus
Allan Hubbard	http://en.wikipedia.org/wiki/Allan_Hubbard_%28Presidential_advisor%29
Allan Lane	http://en.wikipedia.org/wiki/Allan_Lane
Allan Nevins	http://en.wikipedia.org/wiki/Allan_Nevins
Allan Pinkerton	http://en.wikipedia.org/wiki/Allan_Pinkerton
Allard Lowenstein	http://en.wikipedia.org/wiki/Allard_Lowenstein
Allen Boyd	http://en.wikipedia.org/wiki/Allen_Boyd
Allen Drury	http://en.wikipedia.org/wiki/Allen_Drury
Allen Funt	http://en.wikipedia.org/wiki/Allen_Funt
Allen Ginsberg	http://en.wikipedia.org/wiki/Allen_Ginsberg
Allen Hughes	http://en.wikipedia.org/wiki/Allen_Hughes
Allen Iverson	http://en.wikipedia.org/wiki/Allen_Iverson
Allen Klein	http://en.wikipedia.org/wiki/Allen_Klein
Allen Ludden	http://en.wikipedia.org/wiki/Allen_Ludden
Allen Payne	http://en.wikipedia.org/wiki/Allen_Payne
Allen Tate	http://en.wikipedia.org/wiki/Allen_Tate
Allen Toussaint	http://en.wikipedia.org/wiki/Allen_Toussaint
Allen W. Dulles	http://en.wikipedia.org/wiki/Allen_W._Dulles
Allen Weinstein	http://en.wikipedia.org/wiki/Allen_Weinstein
Allison Abbate	http://en.wikipedia.org/wiki/Allison_Abbate
Allison Janney	http://en.wikipedia.org/wiki/Allison_Janney
Allison Mack	http://en.wikipedia.org/wiki/Allison_Mack
Ally Hilfiger	http://en.wikipedia.org/wiki/Ally_Hilfiger
Ally Sheedy	http://en.wikipedia.org/wiki/Ally_Sheedy
Ally Walker	http://en.wikipedia.org/wiki/Ally_Walker
Allyn Joslyn	http://en.wikipedia.org/wiki/Allyn_Joslyn
Allyson Schwartz	http://en.wikipedia.org/wiki/Allyson_Schwartz
Alois Hitler	http://en.wikipedia.org/wiki/Alois_Hitler
Alok Sharma	http://en.wikipedia.org/wiki/Alok_Sharma
Alonso de Castillo Solorzano	http://en.wikipedia.org/wiki/Alonso_de_Castillo_Solorzano
Alonso de Ercilla y Z��iga	http://en.wikipedia.org/wiki/Alonso_de_Ercilla_y_Z%C3%BA%C3%B1iga
Alonzo Mourning	http://en.wikipedia.org/wiki/Alonzo_Mourning
Alphonse Daudet	http://en.wikipedia.org/wiki/Alphonse_Daudet
Alphonse de Lamartine	http://en.wikipedia.org/wiki/Alphonse_de_Lamartine
Alphonso Jackson	http://en.wikipedia.org/wiki/Alphonso_Jackson
Alphonso Taft	http://en.wikipedia.org/wiki/Alphonso_Taft
Althea Flynt	http://en.wikipedia.org/wiki/Althea_Flynt
Althea Gibson	http://en.wikipedia.org/wiki/Althea_Gibson
Alton Brown	http://en.wikipedia.org/wiki/Alton_Brown
Alu Alkhanov	http://en.wikipedia.org/wiki/Alu_Alkhanov
Alun Cairns	http://en.wikipedia.org/wiki/Alun_Cairns
Alun Michael	http://en.wikipedia.org/wiki/Alun_Michael
Alva Myrdal	http://en.wikipedia.org/wiki/Alva_Myrdal
Alvar Aalto	http://en.wikipedia.org/wiki/Alvar_Aalto
�lvaro Colom	http://en.wikipedia.org/wiki/%C1lvaro_Colom
Alvaro Uribe	http://en.wikipedia.org/wiki/Alvaro_Uribe
�lvaro Uribe	http://en.wikipedia.org/wiki/%C1lvaro_Uribe
Alvin Ailey	http://en.wikipedia.org/wiki/Alvin_Ailey
Alvin F. Poussaint	http://en.wikipedia.org/wiki/Alvin_F._Poussaint
Alvin Karpis	http://en.wikipedia.org/wiki/Alvin_Karpis
Alvin Lee	http://en.wikipedia.org/wiki/Alvin_Lee
Alvin Lucier	http://en.wikipedia.org/wiki/Alvin_Lucier
Alvin Toffler	http://en.wikipedia.org/wiki/Alvin_Toffler
Alvin York	http://en.wikipedia.org/wiki/Alvin_York
Alvise Cadamosto	http://en.wikipedia.org/wiki/Alvise_Cadamosto
Alwaleed bin Talal	http://en.wikipedia.org/wiki/Alwaleed_bin_Talal
Aly Khan	http://en.wikipedia.org/wiki/Aly_Khan
Alyson Hannigan	http://en.wikipedia.org/wiki/Alyson_Hannigan
Alyson Michalka	http://en.wikipedia.org/wiki/Alyson_Michalka
Alyssa Milano	http://en.wikipedia.org/wiki/Alyssa_Milano
Amado Nervo	http://en.wikipedia.org/wiki/Amado_Nervo
Amadou Diallo	http://en.wikipedia.org/wiki/Amadou_Diallo
Amadou Toumani Tour�	http://en.wikipedia.org/wiki/Amadou_Toumani_Tour%C3%A9
Amanda Bearse	http://en.wikipedia.org/wiki/Amanda_Bearse
Amanda Blake	http://en.wikipedia.org/wiki/Amanda_Blake
Amanda Bynes	http://en.wikipedia.org/wiki/Amanda_Bynes
Amanda Donohoe	http://en.wikipedia.org/wiki/Amanda_Donohoe
Amanda Pays	http://en.wikipedia.org/wiki/Amanda_Pays
Amanda Peet	http://en.wikipedia.org/wiki/Amanda_Peet
Amanda Plummer	http://en.wikipedia.org/wiki/Amanda_Plummer
Amanda Tapping	http://en.wikipedia.org/wiki/Amanda_Tapping
Amani Abeid Karume	http://en.wikipedia.org/wiki/Amani_Abeid_Karume
Amar Bose	http://en.wikipedia.org/wiki/Amar_Bose
Amartya Sen	http://en.wikipedia.org/wiki/Amartya_Sen
Amazing Kreskin	http://en.wikipedia.org/wiki/Amazing_Kreskin
Amber Benson	http://en.wikipedia.org/wiki/Amber_Benson
Amber Rudd	http://en.wikipedia.org/wiki/Amber_Rudd
Amber Tamblyn	http://en.wikipedia.org/wiki/Amber_Tamblyn
Amber Valletta	http://en.wikipedia.org/wiki/Amber_Valletta
Ambrogio Borgognone	http://en.wikipedia.org/wiki/Ambrogio_Borgognone
Ambroise Par�	http://en.wikipedia.org/wiki/Ambroise_Par%C3%A9
Ambrose Bierce	http://en.wikipedia.org/wiki/Ambrose_Bierce
Ambrose Burnside	http://en.wikipedia.org/wiki/Ambrose_Burnside
Ambrose Philips	http://en.wikipedia.org/wiki/Ambrose_Philips
Amedeo Avogadro	http://en.wikipedia.org/wiki/Amedeo_Avogadro
Amedeo Modigliani	http://en.wikipedia.org/wiki/Amedeo_Modigliani
Amelia Earhart	http://en.wikipedia.org/wiki/Amelia_Earhart
Amelie Mauresmo	http://en.wikipedia.org/wiki/Amelie_Mauresmo
America Ferrera	http://en.wikipedia.org/wiki/America_Ferrera
Amerigo Vespucci	http://en.wikipedia.org/wiki/Amerigo_Vespucci
Amilcare Ponchielli	http://en.wikipedia.org/wiki/Amilcare_Ponchielli
Amin Gemayel	http://en.wikipedia.org/wiki/Amin_Gemayel
Amiri Baraka	http://en.wikipedia.org/wiki/Amiri_Baraka
Amitabh Bachchan	http://en.wikipedia.org/wiki/Amitabh_Bachchan
Ammianus Marcellinus	http://en.wikipedia.org/wiki/Ammianus_Marcellinus
Ammonius Hermiae	http://en.wikipedia.org/wiki/Ammonius_Hermiae
Ammonius Saccas	http://en.wikipedia.org/wiki/Ammonius_Saccas
Amo Houghton	http://en.wikipedia.org/wiki/Amo_Houghton
Amon Goeth	http://en.wikipedia.org/wiki/Amon_Goeth
Amos Rusie	http://en.wikipedia.org/wiki/Amos_Rusie
Amos Tversky	http://en.wikipedia.org/wiki/Amos_Tversky
Amr Mussa	http://en.wikipedia.org/wiki/Amr_Mussa
Amrish Puri	http://en.wikipedia.org/wiki/Amrish_Puri
Amy Acker	http://en.wikipedia.org/wiki/Amy_Acker
Amy Brenneman	http://en.wikipedia.org/wiki/Amy_Brenneman
Amy Carlson	http://en.wikipedia.org/wiki/Amy_Carlson
Amy Carter	http://en.wikipedia.org/wiki/Amy_Carter
Amy Davidson	http://en.wikipedia.org/wiki/Amy_Davidson
Amy Fisher	http://en.wikipedia.org/wiki/Amy_Fisher
Amy Goodman	http://en.wikipedia.org/wiki/Amy_Goodman
Amy Grant	http://en.wikipedia.org/wiki/Amy_Grant
Amy Heckerling	http://en.wikipedia.org/wiki/Amy_Heckerling
Amy Irving	http://en.wikipedia.org/wiki/Amy_Irving
Amy Jacques Garvey	http://en.wikipedia.org/wiki/Amy_Jacques_Garvey
Amy Jo Johnson	http://en.wikipedia.org/wiki/Amy_Jo_Johnson
Amy Klobuchar	http://en.wikipedia.org/wiki/Amy_Klobuchar
Amy Lee	http://en.wikipedia.org/wiki/Amy_Lee
Amy Locane	http://en.wikipedia.org/wiki/Amy_Locane
Amy Lowell	http://en.wikipedia.org/wiki/Amy_Lowell
Amy Madigan	http://en.wikipedia.org/wiki/Amy_Madigan
Amy Pascal	http://en.wikipedia.org/wiki/Amy_Pascal
Amy Pietz	http://en.wikipedia.org/wiki/Amy_Pietz
Amy Poehler	http://en.wikipedia.org/wiki/Amy_Poehler
Amy Ray	http://en.wikipedia.org/wiki/Amy_Ray
Amy Sedaris	http://en.wikipedia.org/wiki/Amy_Sedaris
Amy Smart	http://en.wikipedia.org/wiki/Amy_Smart
Amy Tan	http://en.wikipedia.org/wiki/Amy_Tan
Amy Walter	http://en.wikipedia.org/wiki/Amy_Walters
Amy Winehouse	http://en.wikipedia.org/wiki/Amy_Winehouse
Amy Wynn Pastor	http://en.wikipedia.org/wiki/Amy_Wynn_Pastor
Amy Yasbeck	http://en.wikipedia.org/wiki/Amy_Yasbeck
Ana Hickmann	http://en.wikipedia.org/wiki/Ana_Hickmann
Ana�s Nin	http://en.wikipedia.org/wiki/Ana%C3%AFs_Nin
Anas Sarwar	http://en.wikipedia.org/wiki/Anas_Sarwar
Anastasio Somoza	http://en.wikipedia.org/wiki/Anastasio_Somoza_Debayle
Anatole France	http://en.wikipedia.org/wiki/Anatole_France
Anatole Litvak	http://en.wikipedia.org/wiki/Anatole_Litvak
Anatoli Hrytsenko	http://en.wikipedia.org/wiki/Anatoli_Hrytsenko
Anatoliy Kinakh	http://en.wikipedia.org/wiki/Anatoliy_Kinakh
Anatoly Chubais	http://en.wikipedia.org/wiki/Anatoly_Chubais
Anaximenes of Miletus	http://en.wikipedia.org/wiki/Anaximenes_of_Miletus
Ander Crenshaw	http://en.wikipedia.org/wiki/Ander_Crenshaw
Anders Celsius	http://en.wikipedia.org/wiki/Anders_Celsius
Anders Jonas �ngstr�m	http://en.wikipedia.org/wiki/Anders_Jonas_%C3%85ngstr%C3%B6m
Anderson Cooper	http://en.wikipedia.org/wiki/Anderson_Cooper
Andie MacDowell	http://en.wikipedia.org/wiki/Andie_MacDowell
Andranik Markaryan	http://en.wikipedia.org/wiki/Andranik_Markaryan
Andre 3000	http://en.wikipedia.org/wiki/Andre_3000
Andr� 3000	http://en.wikipedia.org/wiki/Andr%C3%A9_3000
Andr� Aciman	http://en.wikipedia.org/wiki/Andr%C3%A9_Aciman
Andre Agassi	http://en.wikipedia.org/wiki/Andre_Agassi
Andre Braugher	http://en.wikipedia.org/wiki/Andre_Braugher
Andr� Breton	http://en.wikipedia.org/wiki/Andr%C3%A9_Breton
Andr� Carson	http://en.wikipedia.org/wiki/Andr%C3%A9_Carson
Andr� Dacier	http://en.wikipedia.org/wiki/Andr%C3%A9_Dacier
Andr� de Ch�nier	http://en.wikipedia.org/wiki/Andr%C3%A9_de_Ch%C3%A9nier
Andr� Gide	http://en.wikipedia.org/wiki/Andr%C3%A9_Gide
Andr� Malraux	http://en.wikipedia.org/wiki/Andr%C3%A9_Malraux
Andr� Mass�na	http://en.wikipedia.org/wiki/Andr%C3%A9_Mass%C3%A9na
Andr� Maurois	http://en.wikipedia.org/wiki/Andr%C3%A9_Maurois
Andre Norton	http://en.wikipedia.org/wiki/Andre_Norton
Andr� Previn	http://en.wikipedia.org/wiki/Andr%C3%A9_Previn
Andre Soltner	http://en.wikipedia.org/wiki/Andr%C3%A9_Soltner
Andr� the Giant	http://en.wikipedia.org/wiki/Andr%C3%A9_the_Giant
Andr� van Hasselt	http://en.wikipedia.org/wiki/Andr%C3%A9_van_Hasselt
Andrea Barber	http://en.wikipedia.org/wiki/Andrea_Barber
Andrea Bocelli	http://en.wikipedia.org/wiki/Andrea_Bocelli
Andrea Corr	http://en.wikipedia.org/wiki/Andrea_Corr
Andrea del Castagno	http://en.wikipedia.org/wiki/Andrea_del_Castagno
Andrea del Sarto	http://en.wikipedia.org/wiki/Andrea_del_Sarto
Andrea del Verrocchio	http://en.wikipedia.org/wiki/Andrea_del_Verrocchio
Andrea Doria	http://en.wikipedia.org/wiki/Andrea_Doria
Andrea Dworkin	http://en.wikipedia.org/wiki/Andrea_Dworkin
Andrea Jung	http://en.wikipedia.org/wiki/Andrea_Jung
Andrea King	http://en.wikipedia.org/wiki/Andrea_King
Andrea Leadsom	http://en.wikipedia.org/wiki/Andrea_Leadsom
Andrea Mackris	http://en.wikipedia.org/wiki/Andrea_Mackris
Andrea Mantegna	http://en.wikipedia.org/wiki/Andrea_Mantegna
Andrea Martin	http://en.wikipedia.org/wiki/Andrea_Martin
Andrea Mitchell	http://en.wikipedia.org/wiki/Andrea_Mitchell
Andrea Palladio	http://en.wikipedia.org/wiki/Andrea_Palladio
Andrea Parker	http://en.wikipedia.org/wiki/Andrea_Parker
Andrea Pisano	http://en.wikipedia.org/wiki/Andrea_Pisano
Andrea Seabrook	http://en.wikipedia.org/wiki/Andrea_Seabrook
Andrea Yates	http://en.wikipedia.org/wiki/Andrea_Yates
Andreas Hofer	http://en.wikipedia.org/wiki/Andreas_Hofer
Andreas Katsulas	http://en.wikipedia.org/wiki/Andreas_Katsulas
Andreas Osiander	http://en.wikipedia.org/wiki/Andreas_Osiander
Andreas Vesalius	http://en.wikipedia.org/wiki/Andreas_Vesalius
Andr�-Ernest-Modeste Gr�try	http://en.wikipedia.org/wiki/Andr%C3%A9-Ernest-Modeste_Gr%C3%A9try
Andrei Bely	http://en.wikipedia.org/wiki/Andrei_Bely
Andrei Codrescu	http://en.wikipedia.org/wiki/Andrei_Codrescu
Andrei Gromyko	http://en.wikipedia.org/wiki/Andrei_Gromyko
Andrei Sakharov	http://en.wikipedia.org/wiki/Andrei_Sakharov
Andrei Tarkovsky	http://en.wikipedia.org/wiki/Andrei_Tarkovsky
Andr�-Marie Amp�re	http://en.wikipedia.org/wiki/Andr%C3%A9-Marie_Amp%C3%A8re
Andr�s Bello	http://en.wikipedia.org/wiki/Andr%C3%A9s_Bello
Andres Manuel Lopez Obrador	http://en.wikipedia.org/wiki/Andr%C3%A9s_Manuel_L%C3%B3pez_Obrador
Andres Segovia	http://en.wikipedia.org/wiki/Andres_Segovia
Andres Serrano	http://en.wikipedia.org/wiki/Andres_Serrano
Andrew Bell	http://en.wikipedia.org/wiki/Andrew_Bell_%28educationalist%29
Andrew Bingham	http://en.wikipedia.org/wiki/Andrew_Bingham
Andrew Blake	http://en.wikipedia.org/wiki/Andrew_Blake_%28director%29
Andrew Bonar Law	http://en.wikipedia.org/wiki/Andrew_Bonar_Law 
Andrew Bridgen	http://en.wikipedia.org/wiki/Andrew_Bridgen
Andrew Brimmer	http://en.wikipedia.org/wiki/Andrew_Brimmer
Andrew Card	http://en.wikipedia.org/wiki/Andrew_Card
Andrew Carnegie	http://en.wikipedia.org/wiki/Andrew_Carnegie
Andrew Cavendish	http://en.wikipedia.org/wiki/Andrew_Cavendish,_11th_Duke_of_Devonshire
Andrew Cunanan	http://en.wikipedia.org/wiki/Andrew_Cunanan
Andrew Cuomo	http://en.wikipedia.org/wiki/Andrew_Cuomo
Andrew Eldritch	http://en.wikipedia.org/wiki/Andrew_Eldritch
Andrew Fastow	http://en.wikipedia.org/wiki/Andrew_Fastow
Andrew Flintoff	http://en.wikipedia.org/wiki/Andrew_Flintoff
Andrew George	http://en.wikipedia.org/wiki/Andrew_George_%28politician%29
Andrew Gould	http://en.wikipedia.org/wiki/Andrew_Gould
Andrew Griffiths	http://en.wikipedia.org/wiki/Andrew_Griffiths_%28politician%29
Andrew Gwynne	http://en.wikipedia.org/wiki/Andrew_Gwynne
Andrew Heyward	http://en.wikipedia.org/wiki/Andrew_Heyward
Andrew Jackson	http://en.wikipedia.org/wiki/Andrew_Jackson
Andrew Jacobs, Jr.	http://en.wikipedia.org/wiki/Andrew_Jacobs,_Jr.
Andrew Johnson	http://en.wikipedia.org/wiki/Andrew_Johnson
Andrew Jones	http://en.wikipedia.org/wiki/Andrew_Jones_%28politician%29
Andrew Keegan	http://en.wikipedia.org/wiki/Andrew_Keegan
Andrew Lansley	http://en.wikipedia.org/wiki/Andrew_Lansley
Andrew Lawrence	http://en.wikipedia.org/wiki/Andrew_Lawrence_%28actor%29
Andrew Lloyd Webber	http://en.wikipedia.org/wiki/Andrew_Lloyd_Webber
Andrew Marvell	http://en.wikipedia.org/wiki/Andrew_Marvell
Andrew McCarthy	http://en.wikipedia.org/wiki/Andrew_McCarthy
Andrew McKenzie	http://en.wikipedia.org/wiki/Andrew_McKenzie
Andrew Melville	http://en.wikipedia.org/wiki/Andrew_Melville
Andrew Miller	http://en.wikipedia.org/wiki/Andrew_Miller
Andrew Mitchell	http://en.wikipedia.org/wiki/Andrew_Mitchell
Andrew Murrison	http://en.wikipedia.org/wiki/Andrew_Murrison
Andrew Percy	http://en.wikipedia.org/wiki/Andrew_Percy
Andrew Revkin	http://en.wikipedia.org/wiki/Andrew_Revkin
Andrew Reynolds	http://en.wikipedia.org/wiki/Andrew_Reynolds
Andrew Ridgeley	http://en.wikipedia.org/wiki/Andrew_Ridgeley
Andrew Robathan	http://en.wikipedia.org/wiki/Andrew_Robathan
Andrew Roberts	http://en.wikipedia.org/wiki/Andrew_Roberts_%28historian%29
Andrew Rosindell	http://en.wikipedia.org/wiki/Andrew_Rosindell
Andrew Rubin	http://en.wikipedia.org/wiki/Andrew_Rubin
Andrew Selous	http://en.wikipedia.org/wiki/Andrew_Selous
Andrew Shue	http://en.wikipedia.org/wiki/Andrew_Shue
Andrew Smith	http://en.wikipedia.org/wiki/Andrew_Smith_%28politician%29
Andrew Stanton	http://en.wikipedia.org/wiki/Andrew_Stanton
Andrew Stephenson	http://en.wikipedia.org/wiki/Andrew_Stephenson
Andrew Stevens	http://en.wikipedia.org/wiki/Andrew_Stevens
Andrew Stunell	http://en.wikipedia.org/wiki/Andrew_Stunell
Andrew Sullivan	http://en.wikipedia.org/wiki/Andrew_Sullivan
Andrew Tanenbaum	http://en.wikipedia.org/wiki/Andrew_Tanenbaum
Andrew Turner	http://en.wikipedia.org/wiki/Andrew_Turner_%28politician%29
Andrew Tyrie	http://en.wikipedia.org/wiki/Andrew_Tyrie
Andrew V. McLaglen	http://en.wikipedia.org/wiki/Andrew_V._McLaglen
Andrew Vachss	http://en.wikipedia.org/wiki/Andrew_Vachss
Andrew von Eschenbach	http://en.wikipedia.org/wiki/Andrew_von_Eschenbach
Andrew W. Mellon	http://en.wikipedia.org/wiki/Andrew_W._Mellon
Andrew Weil	http://en.wikipedia.org/wiki/Andrew_Weil
Andrew Wiles	http://en.wikipedia.org/wiki/Andrew_Wiles
Andrew Wilson	http://en.wikipedia.org/wiki/Andrew_Wilson_%28actor%29
Andrew Wyeth	http://en.wikipedia.org/wiki/Andrew_Wyeth
Andrew Young	http://en.wikipedia.org/wiki/Andrew_Young
Andrian Nikolayev	http://en.wikipedia.org/wiki/Andrian_Nikolayev
Andrius Kubilius	http://en.wikipedia.org/wiki/Andrius_Kubilius
Andriy Shevchenko	http://en.wikipedia.org/wiki/Andriy_Shevchenko
Andrus Ansip	http://en.wikipedia.org/wiki/Andrus_Ansip
Andy Bell	http://en.wikipedia.org/wiki/Andy_Bell_%28musician%29
Andy Bell	http://en.wikipedia.org/wiki/Andy_Bell_%28singer%29
Andy Burnham	http://en.wikipedia.org/wiki/Andy_Burnham
Andy Devine	http://en.wikipedia.org/wiki/Andy_Devine
Andy Dick	http://en.wikipedia.org/wiki/Andy_Dick
Andy Fairweather-Low	http://en.wikipedia.org/wiki/Andy_Fairweather-Low
Andy Garcia	http://en.wikipedia.org/wiki/Andy_Garcia
Andy Gibb	http://en.wikipedia.org/wiki/Andy_Gibb
Andy Griffith	http://en.wikipedia.org/wiki/Andy_Griffith
Andy Griffiths	http://en.wikipedia.org/wiki/Andy_Griffiths
Andy Grove	http://en.wikipedia.org/wiki/Andy_Grove
Andy Hertzfeld	http://en.wikipedia.org/wiki/Andy_Hertzfeld
Andy Ireland	http://en.wikipedia.org/wiki/Andy_Ireland
Andy Kaufman	http://en.wikipedia.org/wiki/Andy_Kaufman
Andy Love	http://en.wikipedia.org/wiki/Andy_Love
Andy Milonakis	http://en.wikipedia.org/wiki/Andy_Milonakis
Andy Partridge	http://en.wikipedia.org/wiki/Andy_Partridge
Andy Richter	http://en.wikipedia.org/wiki/Andy_Richter
Andy Roddick	http://en.wikipedia.org/wiki/Andy_Roddick
Andy Rooney	http://en.wikipedia.org/wiki/Andy_Rooney
Andy Samberg	http://en.wikipedia.org/wiki/Andy_Samberg
Andy Serkis	http://en.wikipedia.org/wiki/Andy_Serkis
Andy Slaughter	http://en.wikipedia.org/wiki/Andy_Slaughter
Andy Summers	http://en.wikipedia.org/wiki/Andy_Summers
Andy Taylor	http://en.wikipedia.org/wiki/Andy_Taylor_%28guitarist%29
Andy Wachowski	http://en.wikipedia.org/wiki/Andy_Wachowski
Andy Warhol	http://en.wikipedia.org/wiki/Andy_Warhol
Andy Williams	http://en.wikipedia.org/wiki/Andy_Williams
Ang Lee	http://en.wikipedia.org/wiki/Ang_Lee
Angel Cordero	http://en.wikipedia.org/wiki/Angel_Cordero
Angel Tompkins	http://en.wikipedia.org/wiki/Angel_Tompkins
Angela Alioto	http://en.wikipedia.org/wiki/Angela_Alioto
Angela Alvarado	http://en.wikipedia.org/wiki/Angela_Alvarado
Angela Bassett	http://en.wikipedia.org/wiki/Angela_Bassett
Angela C. Smith	http://en.wikipedia.org/wiki/Angela_Christine_Smith
Angela Carter	http://en.wikipedia.org/wiki/Angela_Carter
Angela Cartwright	http://en.wikipedia.org/wiki/Angela_Cartwright
Angela Davis	http://en.wikipedia.org/wiki/Angela_Davis
Angela Eagle	http://en.wikipedia.org/wiki/Angela_Eagle
Angela Georgina Burdett-Coutts	http://en.wikipedia.org/wiki/Angela_Georgina_Burdett-Coutts
Angela Lansbury	http://en.wikipedia.org/wiki/Angela_Lansbury
Angela Merkel	http://en.wikipedia.org/wiki/Angela_Merkel
Angela Watkinson	http://en.wikipedia.org/wiki/Angela_Watkinson
Angelina Jolie	http://en.wikipedia.org/wiki/Angelina_Jolie
Angelo Badalamenti	http://en.wikipedia.org/wiki/Angelo_Badalamenti
Angelo Cardinal Sodano	http://en.wikipedia.org/wiki/Angelo_Cardinal_Sodano
Angelo R. Mozilo	http://en.wikipedia.org/wiki/Angelo_R._Mozilo
Angie Bray	http://en.wikipedia.org/wiki/Angie_Bray
Angie Dickinson	http://en.wikipedia.org/wiki/Angie_Dickinson
Angie Everhart	http://en.wikipedia.org/wiki/Angie_Everhart
Angie Harmon	http://en.wikipedia.org/wiki/Angie_Harmon
Angie Stone	http://en.wikipedia.org/wiki/Angie_Stone
Angus MacNeil	http://en.wikipedia.org/wiki/Angus_MacNeil
Angus Robertson	http://en.wikipedia.org/wiki/Angus_Robertson
Angus Scrimm	http://en.wikipedia.org/wiki/Angus_Scrimm
Angus Wilson	http://en.wikipedia.org/wiki/Angus_Wilson
Angus Young	http://en.wikipedia.org/wiki/Angus_Young
Ani DiFranco	http://en.wikipedia.org/wiki/Ani_DiFranco
An�bal Acevedo-Vil�	http://en.wikipedia.org/wiki/An%C3%ADbal_Acevedo-Vil%C3%A1
An�bal Cavaco Silva	http://en.wikipedia.org/wiki/An%C3%ADbal_Cavaco_Silva
Anil Kapoor	http://en.wikipedia.org/wiki/Anil_Kapoor
Anil Kumble	http://en.wikipedia.org/wiki/Anil_Kumble
Anissa Jones	http://en.wikipedia.org/wiki/Anissa_Jones
Anita Baker	http://en.wikipedia.org/wiki/Anita_Baker
Anita Brookner	http://en.wikipedia.org/wiki/Anita_Brookner
Anita Bryant	http://en.wikipedia.org/wiki/Anita_Bryant
Anita Desai	http://en.wikipedia.org/wiki/Anita_Desai
Anita Ekberg	http://en.wikipedia.org/wiki/Anita_Ekberg
Anita Hill	http://en.wikipedia.org/wiki/Anita_Hill
Anita Loos	http://en.wikipedia.org/wiki/Anita_Loos
Anita O'Day	http://en.wikipedia.org/wiki/Anita_O%27Day
Anita Page	http://en.wikipedia.org/wiki/Anita_Page
Anita Pointer	http://en.wikipedia.org/wiki/Anita_Pointer
Anita W. Addison	http://en.wikipedia.org/wiki/Anita_W._Addison
Anjelica Huston	http://en.wikipedia.org/wiki/Anjelica_Huston
Ann B. Davis	http://en.wikipedia.org/wiki/Ann_B._Davis
Ann Beattie	http://en.wikipedia.org/wiki/Ann_Beattie
Ann Blyth	http://en.wikipedia.org/wiki/Ann_Blyth
Ann Clwyd	http://en.wikipedia.org/wiki/Ann_Clwyd
Ann Coffey	http://en.wikipedia.org/wiki/Ann_Coffey
Ann Coulter	http://en.wikipedia.org/wiki/Ann_Coulter
Ann Curry	http://en.wikipedia.org/wiki/Ann_Curry
Ann Dore McLaughlin	http://en.wikipedia.org/wiki/Ann_Dore_McLaughlin
Ann Druyan	http://en.wikipedia.org/wiki/Ann_Druyan
Ann Jillian	http://en.wikipedia.org/wiki/Ann_Jillian
Ann Kirkpatrick	http://en.wikipedia.org/wiki/Ann_Kirkpatrick
Ann Landers	http://en.wikipedia.org/wiki/Ann_Landers
Ann Magnuson	http://en.wikipedia.org/wiki/Ann_Magnuson
Ann McKechin	http://en.wikipedia.org/wiki/Ann_McKechin
Ann Miller	http://en.wikipedia.org/wiki/Ann_Miller
Ann Petry	http://en.wikipedia.org/wiki/Ann_Petry
Ann Radcliffe	http://en.wikipedia.org/wiki/Ann_Radcliffe
Ann Richards	http://en.wikipedia.org/wiki/Ann_Richards
Ann Robinson	http://en.wikipedia.org/wiki/Ann_Robinson
Ann Rule	http://en.wikipedia.org/wiki/Ann_Rule
Ann Rutherford	http://en.wikipedia.org/wiki/Ann_Rutherford
Ann Sheridan	http://en.wikipedia.org/wiki/Ann_Sheridan
Ann Sothern	http://en.wikipedia.org/wiki/Ann_Sothern
Ann Veneman	http://en.wikipedia.org/wiki/Ann_Veneman
Ann Wedgeworth	http://en.wikipedia.org/wiki/Ann_Wedgeworth
Ann Wilson	http://en.wikipedia.org/wiki/Ann_Wilson
Anna Akhmatova	http://en.wikipedia.org/wiki/Anna_Akhmatova
Anna Chlumsky	http://en.wikipedia.org/wiki/Anna_Chlumsky
Anna Deavere Smith	http://en.wikipedia.org/wiki/Anna_Deavere_Smith
Anna Eshoo	http://en.wikipedia.org/wiki/Anna_Eshoo
Anna Faris	http://en.wikipedia.org/wiki/Anna_Faris
Anna Freud	http://en.wikipedia.org/wiki/Anna_Freud
Anna Friel	http://en.wikipedia.org/wiki/Anna_Friel
Anna Kournikova	http://en.wikipedia.org/wiki/Anna_Kournikova
Anna Lee	http://en.wikipedia.org/wiki/Anna_Lee
Anna Lindh	http://en.wikipedia.org/wiki/Anna_Lindh
Anna Magnani	http://en.wikipedia.org/wiki/Anna_Magnani
Anna Maria Alberghetti	http://en.wikipedia.org/wiki/Anna_Maria_Alberghetti
Anna May Wong	http://en.wikipedia.org/wiki/Anna_May_Wong
Anna Neagle	http://en.wikipedia.org/wiki/Anna_Neagle
Anna Nicole Smith	http://en.wikipedia.org/wiki/Anna_Nicole_Smith
Anna Paquin	http://en.wikipedia.org/wiki/Anna_Paquin
Anna Quindlen	http://en.wikipedia.org/wiki/Anna_Quindlen
Anna Soubry	http://en.wikipedia.org/wiki/Anna_Soubry
Anna Sten	http://en.wikipedia.org/wiki/Anna_Sten
Anna Waronker	http://en.wikipedia.org/wiki/Anna_Waronker
Annabella Sciorra	http://en.wikipedia.org/wiki/Annabella_Sciorra
Annabeth Gish	http://en.wikipedia.org/wiki/Annabeth_Gish
AnnaLee Saxenian	http://en.wikipedia.org/wiki/AnnaLee_Saxenian
Annalise Braakensiek	http://en.wikipedia.org/wiki/Annalise_Braakensiek
Anne Alvaro	http://en.wikipedia.org/wiki/Anne_Alvaro
Anne Archer	http://en.wikipedia.org/wiki/Anne_Archer
Anne Bancroft	http://en.wikipedia.org/wiki/Anne_Bancroft
Anne Baxter	http://en.wikipedia.org/wiki/Anne_Baxter
Anne Begg	http://en.wikipedia.org/wiki/Anne_Begg
Anne Boleyn	http://en.wikipedia.org/wiki/Anne_Boleyn
Anne Boquet	http://en.wikipedia.org/wiki/Anne_Boquet
Anne Bracegirdle	http://en.wikipedia.org/wiki/Anne_Bracegirdle
Anne Bradstreet	http://en.wikipedia.org/wiki/Anne_Bradstreet
Anne Dudley	http://en.wikipedia.org/wiki/Anne_Dudley
Anne Francine	http://en.wikipedia.org/wiki/Anne_Francine
Anne Francis	http://en.wikipedia.org/wiki/Anne_Francis
Anne Frank	http://en.wikipedia.org/wiki/Anne_Frank
Anne Gorsuch	http://en.wikipedia.org/wiki/Anne_Gorsuch
Anne Gwynne	http://en.wikipedia.org/wiki/Anne_Gwynne
Anne Hathaway	http://en.wikipedia.org/wiki/Anne_Hathaway_%28actress%29
Anne Heche	http://en.wikipedia.org/wiki/Anne_Heche
Anne Jeffreys	http://en.wikipedia.org/wiki/Anne_Jeffreys
Anne L. Armstrong	http://en.wikipedia.org/wiki/Anne_L._Armstrong
Anne Lef�vre	http://en.wikipedia.org/wiki/Anne_Lef%C3%A8vre
Anne M. Mulcahy	http://en.wikipedia.org/wiki/Anne_M._Mulcahy
Anne Main	http://en.wikipedia.org/wiki/Anne_Main
Anne McCaffrey	http://en.wikipedia.org/wiki/Anne_McCaffrey
Anne McGuire	http://en.wikipedia.org/wiki/Anne_McGuire
Anne Meara	http://en.wikipedia.org/wiki/Anne_Meara
Anne Milton	http://en.wikipedia.org/wiki/Anne_Milton
Anne Morris	http://en.wikipedia.org/wiki/Anne-Marie_Morris
Anne Morrow Lindbergh	http://en.wikipedia.org/wiki/Anne_Morrow_Lindbergh
Anne Murray	http://en.wikipedia.org/wiki/Anne_Murray
Anne Northup	http://en.wikipedia.org/wiki/Anne_Northup
Anne Oldfield	http://en.wikipedia.org/wiki/Anne_Oldfield
Anne Parrish	http://en.wikipedia.org/wiki/Anne_Parrish
Anne Revere	http://en.wikipedia.org/wiki/Anne_Revere
Anne Rice	http://en.wikipedia.org/wiki/Anne_Rice
Anne Roiphe	http://en.wikipedia.org/wiki/Anne_Roiphe
Anne Sexton	http://en.wikipedia.org/wiki/Anne_Sexton
Anne Shirley	http://en.wikipedia.org/wiki/Anne_Shirley_%28actress%29
Anne Sullivan	http://en.wikipedia.org/wiki/Anne_Sullivan
Anne Tyler	http://en.wikipedia.org/wiki/Anne_Tyler
Anne-Marie Johnson	http://en.wikipedia.org/wiki/Anne-Marie_Johnson
Annette Bening	http://en.wikipedia.org/wiki/Annette_Bening
Annette Brooke	http://en.wikipedia.org/wiki/Annette_Brooke
Annette Dionne	http://en.wikipedia.org/wiki/Annette_Dionne
Annette Funicello	http://en.wikipedia.org/wiki/Annette_Funicello
Annette Lu	http://en.wikipedia.org/wiki/Annette_Lu
Annette O'Toole	http://en.wikipedia.org/wiki/Annette_O%27Toole
Annette Strauss	http://en.wikipedia.org/wiki/Annette_Strauss
Annette Zilinskas	http://en.wikipedia.org/wiki/Annette_Zilinskas
Annie Besant	http://en.wikipedia.org/wiki/Annie_Besant
Annie Dillard	http://en.wikipedia.org/wiki/Annie_Dillard
Annie Leibovitz	http://en.wikipedia.org/wiki/Annie_Leibovitz
Annie Lennox	http://en.wikipedia.org/wiki/Annie_Lennox
Annie Oakley	http://en.wikipedia.org/wiki/Annie_Oakley
Annie Potts	http://en.wikipedia.org/wiki/Annie_Potts
Anni-Frid Lyngstad	http://en.wikipedia.org/wiki/Anni-Frid_Lyngstad
Anote Tong	http://en.wikipedia.org/wiki/Anote_Tong
Anouk Aim�e	http://en.wikipedia.org/wiki/Anouk_Aim%C3%A9e
Anoushka Shankar	http://en.wikipedia.org/wiki/Anoushka_Shankar
Ansel Adams	http://en.wikipedia.org/wiki/Ansel_Adams
Anson Burlingame	http://en.wikipedia.org/wiki/Anson_Burlingame
Anson Williams	http://en.wikipedia.org/wiki/Anson_Williams
Ante Gotovina	http://en.wikipedia.org/wiki/Ante_Gotovina
Anthea Turner	http://en.wikipedia.org/wiki/Anthea_Turner
Anthony � Wood	http://en.wikipedia.org/wiki/Anthony_Wood
Anthony A. Williams	http://en.wikipedia.org/wiki/Anthony_A._Williams
Anthony Anderson	http://en.wikipedia.org/wiki/Anthony_Anderson
Anthony Andrews	http://en.wikipedia.org/wiki/Anthony_Andrews
Anthony Babington	http://en.wikipedia.org/wiki/Anthony_Babington
Anthony Barber	http://en.wikipedia.org/wiki/Anthony_Barber
Anthony Blunt	http://en.wikipedia.org/wiki/Anthony_Blunt
Anthony Bourdain	http://en.wikipedia.org/wiki/Anthony_Bourdain
Anthony Braxton	http://en.wikipedia.org/wiki/Anthony_Braxton
Anthony Burgess	http://en.wikipedia.org/wiki/Anthony_Burgess
Anthony C. Beilenson	http://en.wikipedia.org/wiki/Anthony_C._Beilenson
Anthony Clark	http://en.wikipedia.org/wiki/Anthony_Clark_%28actor%29
Anthony Collins	http://en.wikipedia.org/wiki/Anthony_Collins
Anthony Daniels	http://en.wikipedia.org/wiki/Anthony_Daniels
Anthony Doerr	http://en.wikipedia.org/wiki/Anthony_Doerr
Anthony Eden	http://en.wikipedia.org/wiki/Anthony_Eden
Anthony Edwards	http://en.wikipedia.org/wiki/Anthony_Edwards
Anthony Frederick Augustus Sandys	http://en.wikipedia.org/wiki/Anthony_Frederick_Augustus_Sandys
Anthony Geary	http://en.wikipedia.org/wiki/Anthony_Geary
Anthony Head	http://en.wikipedia.org/wiki/Anthony_Head
Anthony Heald	http://en.wikipedia.org/wiki/Anthony_Heald
Anthony Hecht	http://en.wikipedia.org/wiki/Anthony_Hecht
Anthony Hopkins	http://en.wikipedia.org/wiki/Anthony_Hopkins
Anthony J. Leggett	http://en.wikipedia.org/wiki/Anthony_J._Leggett
Anthony J. Principi	http://en.wikipedia.org/wiki/Anthony_J._Principi
Anthony Kennedy	http://en.wikipedia.org/wiki/Anthony_Kennedy
Anthony Kiedis	http://en.wikipedia.org/wiki/Anthony_Kiedis
Anthony Lake	http://en.wikipedia.org/wiki/Anthony_Lake
Anthony LaPaglia	http://en.wikipedia.org/wiki/Anthony_LaPaglia
Anthony Mann	http://en.wikipedia.org/wiki/Anthony_Mann
Anthony Michael Hall	http://en.wikipedia.org/wiki/Anthony_Michael_Hall
Anthony Minghella	http://en.wikipedia.org/wiki/Anthony_Minghella
Anthony Moore	http://en.wikipedia.org/wiki/Anthony_Moore
Anthony Peeler	http://en.wikipedia.org/wiki/Anthony_Peeler
Anthony Perkins	http://en.wikipedia.org/wiki/Anthony_Perkins
Anthony Powell	http://en.wikipedia.org/wiki/Anthony_Powell
Anthony Quayle	http://en.wikipedia.org/wiki/Anthony_Quayle
Anthony Quinn	http://en.wikipedia.org/wiki/Anthony_Quinn
Anthony Rapp	http://en.wikipedia.org/wiki/Anthony_Rapp
Anthony Romero	http://en.wikipedia.org/wiki/Anthony_Romero
Anthony Russell	http://en.wikipedia.org/wiki/Anthony_Russell
Anthony Shaffer	http://en.wikipedia.org/wiki/Anthony_Shaffer
Anthony Steel	http://en.wikipedia.org/wiki/Anthony_Steel_%28actor%29
Anthony Trollope	http://en.wikipedia.org/wiki/Anthony_Trollope
Anthony Van Dyck	http://en.wikipedia.org/wiki/Anthony_Van_Dyck
Anthony Wayne	http://en.wikipedia.org/wiki/Anthony_Wayne
Anthony Weiner	http://en.wikipedia.org/wiki/Anthony_Weiner
Anthony Zerbe	http://en.wikipedia.org/wiki/Anthony_Zerbe
Anthony Zinni	http://en.wikipedia.org/wiki/Anthony_Zinni
Antoine de Bourbon	http://en.wikipedia.org/wiki/Antoine_de_Bourbon
Antoine de Saint-Exup�ry	http://en.wikipedia.org/wiki/Antoine_de_Saint-Exup%C3%A9ry
Antoine Fran�ois Fourcroy	http://en.wikipedia.org/wiki/Antoine_Fran%C3%A7ois_Fourcroy
Antoine Fuqua	http://en.wikipedia.org/wiki/Antoine_Fuqua
Antoine Watteau	http://en.wikipedia.org/wiki/Antoine_Watteau
Antoine-J�r�me Balard	http://en.wikipedia.org/wiki/Antoine-J%C3%A9r%C3%B4me_Balard
Antoine-Laurent de Lavoisier	http://en.wikipedia.org/wiki/Antoine-Laurent_de_Lavoisier
Antoinette Deshouli�res	http://en.wikipedia.org/wiki/Antoinette_Deshouli%C3%A8res
Anton Bruckner	http://en.wikipedia.org/wiki/Anton_Bruckner
Anton Chekhov	http://en.wikipedia.org/wiki/Anton_Chekhov
Anton LaVey	http://en.wikipedia.org/wiki/Anton_LaVey
Anton Rubinstein	http://en.wikipedia.org/wiki/Anton_Rubinstein
Anton van Leeuwenhoek	http://en.wikipedia.org/wiki/Anton_van_Leeuwenhoek
Anton Webern	http://en.wikipedia.org/wiki/Anton_Webern
Antoni Gaudi	http://en.wikipedia.org/wiki/Antoni_Gaud%C3%AD
Antonin Dvorak	http://en.wikipedia.org/wiki/Anton%C3%ADn_Dvo%C5%99%C3%A1k
Antonin Scalia	ttp://en.wikipedia.org/wiki/Antonin_Scalia
Antonine Maillet	http://en.wikipedia.org/wiki/Antonine_Maillet
Antoninus Pius	http://en.wikipedia.org/wiki/Antoninus_Pius
Antonio Banderas	http://en.wikipedia.org/wiki/Antonio_Banderas
Antonio Canova	http://en.wikipedia.org/wiki/Antonio_Canova
Antonio Carlos Jobim	http://en.wikipedia.org/wiki/Antonio_Carlos_Jobim
Ant�nio de Oliveira Salazar	http://en.wikipedia.org/wiki/Ant%C3%B3nio_de_Oliveira_Salazar
Ant�nio Diniz da Cruz e Silva	http://en.wikipedia.org/wiki/Ant%C3%B3nio_Diniz_da_Cruz_e_Silva
Ant�nio Feliciano de Castilho	http://en.wikipedia.org/wiki/Ant%C3%B3nio_Feliciano_de_Castilho
Antonio Fogazzaro	http://en.wikipedia.org/wiki/Antonio_Fogazzaro
Antonio Genovesi	http://en.wikipedia.org/wiki/Antonio_Genovesi
Antonio Gramsci	http://en.wikipedia.org/wiki/Antonio_Gramsci
Ant�nio Guterres	http://en.wikipedia.org/wiki/Ant%C3%B3nio_Guterres
Antonio Guzm�n Blanco	http://en.wikipedia.org/wiki/Antonio_Guzm%C3%A1n_Blanco
Antonio L�pez de Santa Anna	http://en.wikipedia.org/wiki/Antonio_L%C3%B3pez_de_Santa_Anna
Antonio Machado	http://en.wikipedia.org/wiki/Antonio_Machado
Antonio Moreno	http://en.wikipedia.org/wiki/Antonio_Moreno
Ant�nio �scar Carmona	http://en.wikipedia.org/wiki/Ant%C3%B3nio_%C3%93scar_Carmona
Ant�nio Ramalho Eanes	http://en.wikipedia.org/wiki/Ant%C3%B3nio_Ramalho_Eanes
Antonio Sabato, Jr.	http://en.wikipedia.org/wiki/Antonio_Sabato,_Jr.
Antonio Saca	http://en.wikipedia.org/wiki/Antonio_Saca
Antonio Salieri	http://en.wikipedia.org/wiki/Antonio_Salieri
Antonio Stradivari	http://en.wikipedia.org/wiki/Antonio_Stradivari
Antonio Tabucchi	http://en.wikipedia.org/wiki/Antonio_Tabucchi
Antonio Taguba	http://en.wikipedia.org/wiki/Antonio_Taguba
Antonio Villaraigosa	http://en.wikipedia.org/wiki/Antonio_Villaraigosa
Antonio Vivaldi	http://en.wikipedia.org/wiki/Antonio_Vivaldi
Antony Flew	http://en.wikipedia.org/wiki/Antony_Flew
Antony Hegarty	http://en.wikipedia.org/wiki/Antony_Hegarty
Antony Hewish	http://en.wikipedia.org/wiki/Antony_Hewish
Anushevan Danielian	http://en.wikipedia.org/wiki/Anushavan_Danielyan
Anwar Sadat	http://en.wikipedia.org/wiki/Anwar_Sadat
Anya Seton	http://en.wikipedia.org/wiki/Anya_Seton
Anzia Yezierska	http://en.wikipedia.org/wiki/Anya_Seton
Aphra Behn	http://en.wikipedia.org/wiki/Aphra_Behn
Apisai Ielemia	http://en.wikipedia.org/wiki/Apisai_Ielemia
Apolo Nsibambi	http://en.wikipedia.org/wiki/Apolo_Nsibambi
April Glaspie	http://en.wikipedia.org/wiki/April_Glaspie
Ara Parseghian	http://en.wikipedia.org/wiki/Ara_Parseghian
Arabella Stuart	http://en.wikipedia.org/wiki/Arabella_Stuart
Aram Khachaturian	http://en.wikipedia.org/wiki/Aram_Khachaturian
Arcangelo Corelli	http://en.wikipedia.org/wiki/Arcangelo_Corelli
Archer J. P. Martin	http://en.wikipedia.org/wiki/Archer_John_Porter_Martin
Archibald Campbell Tait	http://en.wikipedia.org/wiki/Archibald_Campbell_Tait
Archibald Cox	http://en.wikipedia.org/wiki/Archibald_Cox
Archibald Johnston	http://en.wikipedia.org/wiki/Archibald_Johnston
Archibald Macleish	http://en.wikipedia.org/wiki/Archibald_Macleish
Archibald Philip Primrose	http://en.wikipedia.org/wiki/Archibald_Philip_Primrose
Archibald Wavell	http://en.wikipedia.org/wiki/Archibald_Wavell
Archie Mayo	http://en.wikipedia.org/wiki/Archie_Mayo
Archie Shepp	http://en.wikipedia.org/wiki/Archie_Shepp
Aretha Franklin	http://en.wikipedia.org/wiki/Aretha_Franklin
Ari Fleischer	http://en.wikipedia.org/wiki/Ari_Fleischer
Arianna Huffington	http://en.wikipedia.org/wiki/Arianna_Huffington
Ariel Durant	http://en.wikipedia.org/wiki/Ariel_Durant
Ariel Sharon	http://en.wikipedia.org/wiki/Ariel_Sharon
Arielle Dombasle	http://en.wikipedia.org/wiki/Arielle_Dombasle
Arielle Tepper	http://en.wikipedia.org/wiki/Arielle_Tepper
Aries Spears	http://en.wikipedia.org/wiki/Aries_Spears
Aristarchus of Samos	http://en.wikipedia.org/wiki/Aristarchus_of_Samos
Aristide Briand	http://en.wikipedia.org/wiki/Aristide_Briand
Aristides Gomes	http://en.wikipedia.org/wiki/Aristides_Gomes
Aristotle Onassis	http://en.wikipedia.org/wiki/Aristotle_Onassis
Arkady Ghoukasyan	http://en.wikipedia.org/wiki/Arkady_Ghoukasyan
Arlan Stangeland	http://en.wikipedia.org/wiki/Arlan_Stangeland
Arlen Specter	http://en.wikipedia.org/wiki/Arlen_Specter
Arlene Dahl	http://en.wikipedia.org/wiki/Arlene_Dahl
Arlene Francis	http://en.wikipedia.org/wiki/Arlene_Francis
Arliss Howard	http://en.wikipedia.org/wiki/Arliss_Howard
Arlo Guthrie	http://en.wikipedia.org/wiki/Arlo_Guthrie
Armand Assante	http://en.wikipedia.org/wiki/Armand_Assante
Armand de Ranc�	http://en.wikipedia.org/wiki/Armand_de_Ranc%C3%A9
Armand Hammer	http://en.wikipedia.org/wiki/Armand_Hammer
Armando Guebuza	http://en.wikipedia.org/wiki/Armando_Guebuza
Armin Meiwes	http://en.wikipedia.org/wiki/Armin_Meiwes
Armin Mueller-Stahl	http://en.wikipedia.org/wiki/Armin_Mueller-Stahl
Armistead Maupin	http://en.wikipedia.org/wiki/Armistead_Maupin
Armstrong Williams	http://en.wikipedia.org/wiki/Armstrong_Williams
Army Archerd	http://en.wikipedia.org/wiki/Army_Archerd
Arna Bontemps	http://en.wikipedia.org/wiki/Arna_Bontemps
Arne Duncan	http://en.wikipedia.org/wiki/Arne_Duncan
Arne Tiselius	http://en.wikipedia.org/wiki/Arne_Tiselius
Arno Penzias	http://en.wikipedia.org/wiki/Arno_Penzias
Arnold Beckman	http://en.wikipedia.org/wiki/Arnold_Beckman
Arnold Bennett	http://en.wikipedia.org/wiki/Arnold_Bennett
Arnold Gingrich	http://en.wikipedia.org/wiki/Arnold_Gingrich
Arnold Newman	http://en.wikipedia.org/wiki/Arnold_Newman
Arnold Palmer	http://en.wikipedia.org/wiki/Arnold_Palmer
Arnold R��tel	http://en.wikipedia.org/wiki/Arnold_R%C3%BC%C3%BCtel
Arnold Schoenberg	http://en.wikipedia.org/wiki/Arnold_Schoenberg
Arnold Schwarzenegger	http://en.wikipedia.org/wiki/Arnold_Schwarzenegger
Arnold Sommerfeld	http://en.wikipedia.org/wiki/Arnold_Sommerfeld
Arnold Toynbee	http://en.wikipedia.org/wiki/Arnold_Toynbee
Arnold Vosloo	http://en.wikipedia.org/wiki/Arnold_Vosloo
Arrigo Boito	http://en.wikipedia.org/wiki/Arrigo_Boito
Arsene Wenger	http://en.wikipedia.org/wiki/Arsene_Wenger
Arsenio Hall	http://en.wikipedia.org/wiki/Arsenio_Hall
Arsenio Martinez Campos	http://en.wikipedia.org/wiki/Arsenio_Martinez_Campos
Art Acord	http://en.wikipedia.org/wiki/Art_Acord
Art Agnos	http://en.wikipedia.org/wiki/Art_Agnos
Art Alexakis	http://en.wikipedia.org/wiki/Art_Alexakis
Art Bell	http://en.wikipedia.org/wiki/Art_Bell
Art Blakey	http://en.wikipedia.org/wiki/Art_Blakey
Art Buchwald	http://en.wikipedia.org/wiki/Art_Buchwald
Art Carney	http://en.wikipedia.org/wiki/Art_Carney
Art Donovan	http://en.wikipedia.org/wiki/Art_Donovan
Art Fleming	http://en.wikipedia.org/wiki/Art_Fleming
Art Garfunkel	http://en.wikipedia.org/wiki/Art_Garfunkel
Art James	http://en.wikipedia.org/wiki/Art_Jamesn
Art Linkletter	http://en.wikipedia.org/wiki/Art_Linkletter
Art Modell	http://en.wikipedia.org/wiki/Art_Modell
Art Neville	http://en.wikipedia.org/wiki/Art_Neville
Art Rooney	http://en.wikipedia.org/wiki/Art_Rooney
Art Spiegelman	http://en.wikipedia.org/wiki/Art_Spiegelman
Arte Johnson	http://en.wikipedia.org/wiki/Arte_Johnson
Artemas Ward	http://en.wikipedia.org/wiki/Artemas_Ward
Artemisia Gentileschi	http://en.wikipedia.org/wiki/Artemisia_Gentileschi
Artemus Ward	http://en.wikipedia.org/wiki/Artemus_Ward
Arthur "Doc" Barker	http://en.wikipedia.org/wiki/Arthur_Barker
Arthur Agatston	http://en.wikipedia.org/wiki/Arthur_Agatston
Arthur Alexander	http://en.wikipedia.org/wiki/Arthur_Alexander
Arthur Ashe	http://en.wikipedia.org/wiki/Arthur_Ashe
Arthur Askey	http://en.wikipedia.org/wiki/Arthur_Askey
Arthur B. Laffer	http://en.wikipedia.org/wiki/Arthur_B._Laffer
Arthur Balfour	http://en.wikipedia.org/wiki/Arthur_Balfour
Arthur Blank	http://en.wikipedia.org/wiki/Arthur_Blank
Arthur Bremer	http://en.wikipedia.org/wiki/Arthur_Bremer
Arthur Brown	http://en.wikipedia.org/wiki/Arthur_Brown_%28musician%29
Arthur Bryant	http://en.wikipedia.org/wiki/Arthur_Bryant
Arthur C. Clarke	http://en.wikipedia.org/wiki/Arthur_C._Clarke
Arthur C. Nielsen	http://en.wikipedia.org/wiki/Arthur_C._Nielsen
Arthur Conan Doyle	http://en.wikipedia.org/wiki/Arthur_Conan_Doyle
Arthur Conley	http://en.wikipedia.org/wiki/Arthur_Conley
Arthur Dion Hanna	http://en.wikipedia.org/wiki/Arthur_Dion_Hanna
Arthur Dyer Tripp III	http://en.wikipedia.org/wiki/Art_Tripp
Arthur Edward Waite	http://en.wikipedia.org/wiki/Arthur_Edward_Waite
Arthur Fiedler	http://en.wikipedia.org/wiki/Arthur_Fiedler
Arthur Franz	http://en.wikipedia.org/wiki/Arthur_Franz
Arthur Freed	http://en.wikipedia.org/wiki/Arthur_Freed
Arthur Gary Bishop	http://en.wikipedia.org/wiki/Arthur_Gary_Bishop
Arthur Godfrey	http://en.wikipedia.org/wiki/Arthur_Godfrey
Arthur H. Compton	http://en.wikipedia.org/wiki/Arthur_H._Compton
Arthur Hailey	http://en.wikipedia.org/wiki/Arthur_Hailey
Arthur Harden	http://en.wikipedia.org/wiki/Arthur_Harden
Arthur Hayes Sulzberger	http://en.wikipedia.org/wiki/Arthur_Hayes_Sulzberger
Arthur Henderson	http://en.wikipedia.org/wiki/Arthur_Henderson
Arthur Hill	http://en.wikipedia.org/wiki/Arthur_Hill_%28actor%29
Arthur Hiller	http://en.wikipedia.org/wiki/Arthur_Hiller
Arthur Honegger	http://en.wikipedia.org/wiki/Arthur_Honegger
Arthur J. Goldberg	http://en.wikipedia.org/wiki/Arthur_J._Goldberg
Arthur Kennedy	http://en.wikipedia.org/wiki/Arthur_Kennedy_%28actor%29
Arthur Koestler	http://en.wikipedia.org/wiki/Arthur_Koestler
Arthur Kopit	http://en.wikipedia.org/wiki/Arthur_Kopit
Arthur L. Schawlow	http://en.wikipedia.org/wiki/Arthur_L._Schawlow
Arthur Laurents	http://en.wikipedia.org/wiki/Arthur_Laurents
Arthur Levitt	http://en.wikipedia.org/wiki/Arthur_Levitt
Arthur Lowe	http://en.wikipedia.org/wiki/Arthur_Lowe
Arthur Lubin	http://en.wikipedia.org/wiki/Arthur_Lubin
Arthur M. Schlesinger	http://en.wikipedia.org/wiki/Arthur_M._Schlesinger
Arthur Machen	http://en.wikipedia.org/wiki/Arthur_Schlesinger,_Jr.
Arthur Malet	http://en.wikipedia.org/wiki/Arthur_Malet
Arthur Meighen	http://en.wikipedia.org/wiki/Arthur_Meighen
Arthur Miller	http://en.wikipedia.org/wiki/Arthur_Miller
Arthur Murray	http://en.wikipedia.org/wiki/Arthur_Murray
Arthur O. Lovejoy	http://en.wikipedia.org/wiki/Arthur_O._Lovejoy
Arthur Penn	http://en.wikipedia.org/wiki/Arthur_Penn
Arthur Rackham	http://en.wikipedia.org/wiki/Arthur_Rackham
Arthur Rimbaud	http://en.wikipedia.org/wiki/Arthur_Rimbaud
Arthur Rock	http://en.wikipedia.org/wiki/Arthur_Rock
Arthur Schnitzler	http://en.wikipedia.org/wiki/Arthur_Schnitzler
Arthur Schopenhauer	http://en.wikipedia.org/wiki/Arthur_Schopenhauer
Arthur Seyss-Inquart	http://en.wikipedia.org/wiki/Arthur_Seyss-Inquart
Arthur Shawcross	http://en.wikipedia.org/wiki/Arthur_Shawcross
Arthur Sullivan	http://en.wikipedia.org/wiki/Arthur_Sullivan
Arthur Sulzberger, Jr.	http://en.wikipedia.org/wiki/Arthur_Sulzberger,_Jr.
Arthur Symons	http://en.wikipedia.org/wiki/Arthur_Symons
Arthur Treacher	http://en.wikipedia.org/wiki/Treacher
Arthur Vandenberg	http://en.wikipedia.org/wiki/Arthur_Vandenberg
Arthur Wellesley	http://en.wikipedia.org/wiki/Arthur_Wellesley,_1st_Duke_of_Wellington
Arthur Wing Pinero	http://en.wikipedia.org/wiki/Arthur_Wing_Pinero
Arthur Zimmermann	http://en.wikipedia.org/wiki/Arthur_Zimmermann
Artie Lange	http://en.wikipedia.org/wiki/Artie_Lange
Artie Mitchell	http://en.wikipedia.org/wiki/Artie_Mitchell
Artie Shaw	http://en.wikipedia.org/wiki/Artie_Shaw
Arto Lindsay	http://en.wikipedia.org/wiki/Arto_Lindsay
Artturi Virtanen	http://en.wikipedia.org/wiki/Artturi_Virtanen
Artur Axmann	http://en.wikipedia.org/wiki/Artur_Axmann
Artur Davis	http://en.wikipedia.org/wiki/Artur_Davis
Artur Rasizade	http://en.wikipedia.org/wiki/Artur_Rasizade
Artur Rubinstein	http://en.wikipedia.org/wiki/Artur_Rubinstein
Artur Schnabel	http://en.wikipedia.org/wiki/Artur_Schnabel
Arturo Toscanini	http://en.wikipedia.org/wiki/Arturo_Toscanini
Arundhati Roy	http://en.wikipedia.org/wiki/Arundhati_Roy
Ary Barroso	http://en.wikipedia.org/wiki/Ary_Barroso
Asa Gray	http://en.wikipedia.org/wiki/Asa_Gray
Asa Hutchinson	http://en.wikipedia.org/wiki/Asa_Hutchinson
Ashlee Simpson	http://en.wikipedia.org/wiki/Ashlee_Simpson
Ashleigh Banfield	http://en.wikipedia.org/wiki/Ashleigh_Banfield
Ashleigh Brilliant	http://en.wikipedia.org/wiki/Ashleigh_Brilliant
Ashley Harkleroad	http://en.wikipedia.org/wiki/Ashley_Harkleroad
Ashley Judd	http://en.wikipedia.org/wiki/Ashley_Judd
Ashley Montagu	http://en.wikipedia.org/wiki/Ashley_Montagu
Ashley Olsen	http://en.wikipedia.org/wiki/Ashley_Olsen
Ashley Parker Angel	http://en.wikipedia.org/wiki/Ashley_Parker_Angel
Ashley Scott	http://en.wikipedia.org/wiki/Ashley_Scott
Ashley Tisdale	http://en.wikipedia.org/wiki/Ashley_Tisdale
Ashton Kutcher	http://en.wikipedia.org/wiki/Ashton_Kutcher
Asia Argento	http://en.wikipedia.org/wiki/Asia_Argento
Asia Carrera	http://en.wikipedia.org/wiki/Asia_Carrera
Asif Ali Zardari	http://en.wikipedia.org/wiki/Asif_Ali_Zardari
Askar Akayev	http://en.wikipedia.org/wiki/Asif_Ali_Zardari
Atal Bihari Vajpayee	http://en.wikipedia.org/wiki/Atal_Bihari_Vajpayee
Athanasius Kircher	http://en.wikipedia.org/wiki/Athanasius_Kircher
Athina Onassis Roussel	http://en.wikipedia.org/wiki/Athina_Onassis_Roussel
Athol Fugard	http://en.wikipedia.org/wiki/Athol_Fugard
Atom Egoyan	http://en.wikipedia.org/wiki/Atom_Egoyan
Attila the Hun	http://en.wikipedia.org/wiki/Attila_the_Hun
Auberon Waugh	http://en.wikipedia.org/wiki/Auberon_Waugh
Aubrey Beardsley	http://en.wikipedia.org/wiki/Aubrey_Beardsley
Audie England	http://en.wikipedia.org/wiki/Audie_England
Audie Murphy	http://en.wikipedia.org/wiki/Audie_Murphy
Audra Lindley	http://en.wikipedia.org/wiki/Audra_Lindley
Audre Lorde	http://en.wikipedia.org/wiki/Audre_Lorde
Audrey Hepburn	http://en.wikipedia.org/wiki/Audrey_Hepburn
Audrey Landers	http://en.wikipedia.org/wiki/Audrey_Landers
Audrey Meadows	http://en.wikipedia.org/wiki/Audrey_Meadows
Audrey Santo	http://en.wikipedia.org/wiki/Audrey_Santo
Audrey Tautou	http://en.wikipedia.org/wiki/Audrey_Tautou
August Kleinzahler	http://en.wikipedia.org/wiki/August_Kleinzahler
August Strindberg	http://en.wikipedia.org/wiki/August_Strindberg
August Weismann	http://en.wikipedia.org/wiki/August_Weismann
August Wilhelm von Hofmann	http://en.wikipedia.org/wiki/August_Wilhelm_von_Hofmann
August Wilhelm von Schlegel	http://en.wikipedia.org/wiki/August_Wilhelm_von_Schlegel
August Wilson	http://en.wikipedia.org/wiki/August_Wilson
Augusta, Lady Gregory	http://en.wikipedia.org/wiki/Augusta,_Lady_Gregory
Auguste Beernaert	http://en.wikipedia.org/wiki/Auguste_Beernaert
Auguste Comte	http://en.wikipedia.org/wiki/Auguste_Comte
Auguste Escoffier	http://en.wikipedia.org/wiki/Auguste_Escoffier
Auguste Renoir	http://en.wikipedia.org/wiki/Auguste_Renoir
Auguste Rodin	http://en.wikipedia.org/wiki/Auguste_Rodin
Augusten Burroughs	http://en.wikipedia.org/wiki/Augusten_Burroughs
Augustin-Jean Fresnel	http://en.wikipedia.org/wiki/Augustin-Jean_Fresnel
Augustin-Louis Cauchy	http://en.wikipedia.org/wiki/Augustin-Louis_Cauchy
Augusto Pinochet	http://en.wikipedia.org/wiki/Augusto_Pinochet
Augustus Baldwin Longstreet	http://en.wikipedia.org/wiki/Augustus_Baldwin_Longstreet
Augustus De Morgan	http://en.wikipedia.org/wiki/Augustus_De_Morgan
Augustus Egg	http://en.wikipedia.org/wiki/Augustus_Egg
Augustus F. Hawkins	http://en.wikipedia.org/wiki/Augustus_F._Hawkins
Augustus I	http://en.wikipedia.org/wiki/Augustus_I
Augustus II	http://en.wikipedia.org/wiki/Augustus_II_the_Strong
Augustus III	http://en.wikipedia.org/wiki/Augustus_III_of_Poland
Augustus Saint-Gaudens	http://en.wikipedia.org/wiki/Augustus_Saint-Gaudens
Augustus Welby Pugin	http://en.wikipedia.org/wiki/Augustus_Welby_Pugin
Aung San Suu Kyi	http://en.wikipedia.org/wiki/Aung_San_Suu_Kyi
Aurelie Claudel	http://en.wikipedia.org/wiki/Aurelie_Claudel
Austen Chamberlain	http://en.wikipedia.org/wiki/Austen_Chamberlain
Austin J. Murphy	http://en.wikipedia.org/wiki/Austin_J._Murphy
Austin Mitchell	http://en.wikipedia.org/wiki/Austin_Mitchell
Ava Gardner	http://en.wikipedia.org/wiki/Ava_Gardner
Avery Brooks	http://en.wikipedia.org/wiki/Avery_Brooks
Avery Brundage	http://en.wikipedia.org/wiki/Avery_Brundage
Avril Lavigne	http://en.wikipedia.org/wiki/Avril_Lavigne
Axl Rose	http://en.wikipedia.org/wiki/Axl_Rose
Ayatollah Khamenei	http://en.wikipedia.org/wiki/Ayatollah_Khamenei
Ayi Kwei Armah	http://en.wikipedia.org/wiki/Ayi_Kwei_Armah
Aylmer Maude	http://en.wikipedia.org/wiki/Aylmer_Maude
Ayman al-Zawahiri	http://en.wikipedia.org/wiki/Ayman_al-Zawahiri
Ayn Rand	http://en.wikipedia.org/wiki/Ayn_Rand
Aynsley Dunbar	http://en.wikipedia.org/wiki/Aynsley_Dunbar
Ayrton Senna	http://en.wikipedia.org/wiki/Ayrton_Senna
Azali Assoumani	http://en.wikipedia.org/wiki/Azali_Assoumani
Azita Youssefi	http://en.wikipedia.org/wiki/Azita_Youssefi
B. B. King	http://en.wikipedia.org/wiki/B._B._King
B. Carroll Reece	http://en.wikipedia.org/wiki/B._Carroll_Reece
B. D. Wong	http://en.wikipedia.org/wiki/B._D._Wong
B. F. Skinner	http://en.wikipedia.org/wiki/B._F._Skinner
B. J. Habibie	http://en.wikipedia.org/wiki/B._J._Habibie
Babe Ruth	http://en.wikipedia.org/wiki/Babe_Ruth
Babe Zaharias	http://en.wikipedia.org/wiki/Babe_Zaharias
Babrak Karmal	http://en.wikipedia.org/wiki/Babrak_Karmal
Baby Bash	http://en.wikipedia.org/wiki/Baby_Bash
Baby Huey	http://en.wikipedia.org/wiki/Baby_Huey
Baghdadi Mahmudi	http://en.wikipedia.org/wiki/Baghdadi_Mahmudi
Bai Ling	http://en.wikipedia.org/wiki/Bai_Ling
Bainbridge Colby	http://en.wikipedia.org/wiki/Bainbridge_Colby
Bajram Kosumi	http://en.wikipedia.org/wiki/Bajram_Kosumi
Baldassare Castiglione	http://en.wikipedia.org/wiki/Baldassare_Castiglione
Baldassare Galuppi	http://en.wikipedia.org/wiki/Baldassare_Galuppi
Baldassarre Peruzzi	http://en.wikipedia.org/wiki/Baldassarre_Peruzzi
Baldur von Schirach	http://en.wikipedia.org/wiki/Baldur_von_Schirach
Baldwin Spencer	http://en.wikipedia.org/wiki/Baldwin_Spencer
Balfour Stewart	http://en.wikipedia.org/wiki/Balfour_Stewart
Balthazar Getty	http://en.wikipedia.org/wiki/Balthazar_Getty
Bam Margera	http://en.wikipedia.org/wiki/Bam_Margera
Bamir Topi	http://en.wikipedia.org/wiki/Bamir_Topi
Bankim Chandra Chatterji	http://en.wikipedia.org/wiki/Bankim_Chandra_Chatterji
Barack Obama	http://en.wikipedia.org/wiki/Barack_Obama
Barbara A. Mikulski	http://en.wikipedia.org/wiki/Barbara_A._Mikulski
Barbara Amiel	http://en.wikipedia.org/wiki/Barbara_Amiel
Barbara B. Kennelly	http://en.wikipedia.org/wiki/Barbara_B._Kennelly
Barbara Bach	http://en.wikipedia.org/wiki/Barbara_Bach
Barbara Bain	http://en.wikipedia.org/wiki/Barbara_Bain
Barbara Bates	Phttp://en.wikipedia.org/wiki/Barbara_Bates
Barbara Bel Geddes	http://en.wikipedia.org/wiki/Barbara_Bel_Geddes
Barbara Billingsley	http://en.wikipedia.org/wiki/Barbara_Billingsley
Barbara Boxer	http://en.wikipedia.org/wiki/Barbara_Boxer
Barbara Britton	http://en.wikipedia.org/wiki/Barbara_Britton
Barbara Bush	http://en.wikipedia.org/wiki/Barbara_Bush
Barbara Bush	http://en.wikipedia.org/wiki/Barbara_Pierce_Bush
Barbara Carrera	http://en.wikipedia.org/wiki/Barbara_Carrera
Barbara Cartland	http://en.wikipedia.org/wiki/Barbara_Cartland
Barbara Cook	http://en.wikipedia.org/wiki/Barbara_Cook
Barbara Cubin	http://en.wikipedia.org/wiki/Barbara_Cubin
Barbara Eden	http://en.wikipedia.org/wiki/Barbara_Eden
Barbara Ehrenreich	http://en.wikipedia.org/wiki/Barbara_Ehrenreich
Barbara F. Vucanovich	http://en.wikipedia.org/wiki/Barbara_F._Vucanovich
Barbara Feldon	http://en.wikipedia.org/wiki/Barbara_Feldon
Barbara Gaskin	http://en.wikipedia.org/wiki/Barbara_Gaskin
Barbara Hackman Franklin	http://en.wikipedia.org/wiki/Barbara_Hackman_Franklin
Barbara Hale	http://en.wikipedia.org/wiki/Barbara_Hale
Barbara Harris	http://en.wikipedia.org/wiki/Barbara_Harris_%28actress%29
Barbara Hepworth	http://en.wikipedia.org/wiki/Barbara_Hepworth
Barbara Hershey	http://en.wikipedia.org/wiki/Barbara_Hershey
Barbara Jo Allen	http://en.wikipedia.org/wiki/Barbara_Jo_Allen
Barbara Jordan	http://en.wikipedia.org/wiki/Barbara_Jordan
Barbara Keeley	http://en.wikipedia.org/wiki/Barbara_Keeley
Barbara Kent	http://en.wikipedia.org/wiki/Barbara_Kent
Barbara Kingsolver	http://en.wikipedia.org/wiki/Barbara_Kingsolver
Barbara Lee	http://en.wikipedia.org/wiki/Barbara_Lee
Barbara Leigh	http://en.wikipedia.org/wiki/Barbara_Leigh
Barbara Mandrell	http://en.wikipedia.org/wiki/Barbara_Mandrell
Barbara McClintock	http://en.wikipedia.org/wiki/Barbara_McClintock
Barbara Mikulski	http://en.wikipedia.org/wiki/Barbara_Mikulski
Barbara Nichols	http://en.wikipedia.org/wiki/Barbara_Nichols
Barbara Olson	http://en.wikipedia.org/wiki/Barbara_Olson
Barbara O'Neil	http://en.wikipedia.org/wiki/Barbara_O%27Neil
Barbara Parkins	http://en.wikipedia.org/wiki/Barbara_Parkins
Barbara Payton	http://en.wikipedia.org/wiki/Barbara_Payton
Barbara Pym	http://en.wikipedia.org/wiki/Barbara_Pym
Barbara Rush	http://en.wikipedia.org/wiki/Barbara_Rush
Barbara Stanwyck	http://en.wikipedia.org/wiki/Barbara_Stanwyck
Barbara Steele	http://en.wikipedia.org/wiki/Barbara_Steele
Barbara Taylor Bradford	http://en.wikipedia.org/wiki/Barbara_Taylor_Bradford
Barbara Tuchman	http://en.wikipedia.org/wiki/Barbara_Tuchman
Barbara Walters	http://en.wikipedia.org/wiki/Barbara_Walters
Barbara Windsor	http://en.wikipedia.org/wiki/Barbara_Windsor
Barber Conable	http://en.wikipedia.org/wiki/Barber_Conable
Barbet Schroeder	http://en.wikipedia.org/wiki/Barbet_Schroeder
Barbi Benton	http://en.wikipedia.org/wiki/Barbi_Benton
Barbra Streisand	http://en.wikipedia.org/wiki/Barbra_Streisand
Barnabas Sibusiso Dlamini	http://en.wikipedia.org/wiki/Barnabas_Sibusiso_Dlamini
Barnard Hughes	http://en.wikipedia.org/wiki/Barnard_Hughes
Barnett Newman	http://en.wikipedia.org/wiki/Barnett_Newman
Barney Frank	http://en.wikipedia.org/wiki/Barney_Frank
Barney Kessel	http://en.wikipedia.org/wiki/Barney_Kessel
Barney Martin	http://en.wikipedia.org/wiki/Barney_Martin
Barney Oliver	http://en.wikipedia.org/wiki/Barney_Oliver
Baron Hill	http://en.wikipedia.org/wiki/Baron_Hill
Barret Oliver	http://en.wikipedia.org/wiki/Barret_Oliver
Barret Robbins	http://en.wikipedia.org/wiki/Barret_Robbins
Barrett Strong	http://en.wikipedia.org/wiki/Barrett_Strong
Barrington Levy	http://en.wikipedia.org/wiki/Barrington_Levy
Barron Hilton	http://en.wikipedia.org/wiki/Barron_Hilton
Barry Bonds	http://en.wikipedia.org/wiki/Barry_Bonds
Barry Bostwick	http://en.wikipedia.org/wiki/Barry_Bostwick
Barry Commoner	http://en.wikipedia.org/wiki/Barry_Commoner
Barry Corbin	http://en.wikipedia.org/wiki/Barry_Corbin
Barry Davies	http://en.wikipedia.org/wiki/Barry_Davies
Barry Diller	http://en.wikipedia.org/wiki/Barry_Diller
Barry Fitzgerald	http://en.wikipedia.org/wiki/Barry_Fitzgerald
Barry Gardiner	http://en.wikipedia.org/wiki/Barry_Gardiner
Barry Gibb	http://en.wikipedia.org/wiki/Barry_Gibb
Barry Goldwater	http://en.wikipedia.org/wiki/Barry_Goldwater
Barry Guy	http://en.wikipedia.org/wiki/Barry_Guy
Barry Hannah	http://en.wikipedia.org/wiki/Barry_Hannah
Barry Humphries	http://en.wikipedia.org/wiki/Barry_Humphries
Barry Levinson	http://en.wikipedia.org/wiki/Barry_Levinson
Barry Lopez	http://en.wikipedia.org/wiki/Barry_Lopez
Barry Lynn	http://en.wikipedia.org/wiki/Barry_W._Lynn
Barry Manilow	http://en.wikipedia.org/wiki/Barry_Manilow
Barry Mann	http://en.wikipedia.org/wiki/Barry_Mann
Barry McCaffrey	http://en.wikipedia.org/wiki/Barry_McCaffrey
Barry Morse	http://en.wikipedia.org/wiki/Barry_Morse
Barry Nelson	http://en.wikipedia.org/wiki/Barry_Nelson
Barry Pepper	http://en.wikipedia.org/wiki/Barry_Pepper
Barry Sanders	http://en.wikipedia.org/wiki/Barry_Sanders
Barry Sheerman	http://en.wikipedia.org/wiki/Barry_Sheerman
Barry Sonnenfeld	http://en.wikipedia.org/wiki/Barry_Sonnenfeld
Barry Sullivan	http://en.wikipedia.org/wiki/Barry_Sullivan_%28actor%29
Barry Switzer	http://en.wikipedia.org/wiki/Barry_Switzer
Barry Unsworth	http://en.wikipedia.org/wiki/Barry_Unsworth
Barry Van Dyke	http://en.wikipedia.org/wiki/Barry_Van_Dyke
Barry Watson	http://en.wikipedia.org/wiki/Barry_Watson_%28actor%29
Barry White	http://en.wikipedia.org/wiki/Barry_White
Barry Williams	http://en.wikipedia.org/wiki/Barry_Williams
Barry Wood	http://en.wikipedia.org/wiki/Barry_Wood_%28interior_designer%29
Barry Zito	http://en.wikipedia.org/wiki/Barry_Zito
Bart Braverman	http://en.wikipedia.org/wiki/Bart_Braverman
Bart Freundlich	http://en.wikipedia.org/wiki/Bart_Freundlich
Bart Giamatti	http://en.wikipedia.org/wiki/Bart_Giamatti
Bart Gordon	http://en.wikipedia.org/wiki/Bart_Gordon
Bart Starr	http://en.wikipedia.org/wiki/Bart_Starr
Bart Stupak	http://en.wikipedia.org/wiki/Bart_Stupak
Barth�lemy-Prosper Enfantin	http://en.wikipedia.org/wiki/Barth%C3%A9lemy-Prosper_Enfantin
Bartholomew Diaz	http://en.wikipedia.org/wiki/Bartholomew_Diaz
Bartholomew I	http://en.wikipedia.org/wiki/Bartholomew_I
Bartolom� Esteban Murillo	http://en.wikipedia.org/wiki/Bartolom%C3%A9_Esteban_Murillo
Bartolommeo Ammannati	http://en.wikipedia.org/wiki/Bartolommeo_Ammannati
Baruch de Spinoza	http://en.wikipedia.org/wiki/Baruch_de_Spinoza
Bashar al-Assad	http://en.wikipedia.org/wiki/Bashar_al-Assad
Basil Dearden	http://en.wikipedia.org/wiki/Basil_Dearden
Basil King	http://en.wikipedia.org/wiki/Basil_King
Basil Liddell Hart	http://en.wikipedia.org/wiki/Basil_Liddell_Hart
Basil Rathbone	http://en.wikipedia.org/wiki/Basil_Rathbone
Baudouin I	http://en.wikipedia.org/wiki/Baudouin_I
Bay Buchanan	http://en.wikipedia.org/wiki/Bay_Buchanan
Bayard Rustin	http://en.wikipedia.org/wiki/Bayard_Rustin
Bayard Taylor	http://en.wikipedia.org/wiki/Bayard_Taylor
Bayezid I	http://en.wikipedia.org/wiki/Bayezid_I
Bayezid II	http://en.wikipedia.org/wiki/Bayezid_II
Baz Luhrmann	http://en.wikipedia.org/wiki/Baz_Luhrmann
Bea Arthur	http://en.wikipedia.org/wiki/Bea_Arthur
Bea Benaderet	http://en.wikipedia.org/wiki/Bea_Benaderet
Beanie Sigel	http://en.wikipedia.org/wiki/Beanie_Sigel
Bear Bryant	http://en.wikipedia.org/wiki/Bear_Bryant
Beatrice Cenci	http://en.wikipedia.org/wiki/Beatrice_Cenci
Beatrice Straight	http://en.wikipedia.org/wiki/Beatrice_Straight
Beatrice Wood	http://en.wikipedia.org/wiki/Beatrice_Wood
Beatrix of the Netherlands	http://en.wikipedia.org/wiki/Beatrix_of_the_Netherlands
Beatrix Potter	http://en.wikipedia.org/wiki/Beatrix_Potter
Beau Boulter	http://en.wikipedia.org/wiki/Beau_Boulter
Beau Bridges	http://en.wikipedia.org/wiki/Beau_Bridges
Beau Brummell	http://en.wikipedia.org/wiki/Beau_Brummell
Bebe Buell	http://en.wikipedia.org/wiki/Bebe_Buell
Bebe Daniels	http://en.wikipedia.org/wiki/Bebe_Daniels
Bebe Neuwirth	http://en.wikipedia.org/wiki/Bebe_Neuwirth
Bec Cartwright	http://en.wikipedia.org/wiki/Bec_Cartwright
Bedrich Smetana	http://en.wikipedia.org/wiki/Bedrich_Smetana
Beenie Man	http://en.wikipedia.org/wiki/Beenie_Man
Bei Dao	http://en.wikipedia.org/wiki/Bei_Dao
Bela Bartok	http://en.wikipedia.org/wiki/Bela_Bartok
Bela Fleck	http://en.wikipedia.org/wiki/Bela_Fleck
Bela Lugosi	http://en.wikipedia.org/wiki/Bela_Lugosi
Belinda Carlisle	http://en.wikipedia.org/wiki/Belinda_Carlisle
Belinda Lee	http://en.wikipedia.org/wiki/Belinda_Lee
bell hooks	http://en.wikipedia.org/wiki/bell_hooks
Ben Affleck	http://en.wikipedia.org/wiki/Ben_Affleck
Ben Bernanke	http://en.wikipedia.org/wiki/Ben_Bernanke
Ben Blaz	http://en.wikipedia.org/wiki/Ben_Blaz
Ben Bova	http://en.wikipedia.org/wiki/Ben_Bova
Ben Bradlee	http://en.wikipedia.org/wiki/Ben_Bradlee
Ben Bradshaw	http://en.wikipedia.org/wiki/Ben_Bradshaw
Ben Browder	http://en.wikipedia.org/wiki/Ben_Browder
Ben Cardin	http://en.wikipedia.org/wiki/Ben_Cardin
Ben Chandler	http://en.wikipedia.org/wiki/Ben_Chandler
Ben Chaplin	http://en.wikipedia.org/wiki/Ben_Chaplin
Ben Cohen	http://en.wikipedia.org/wiki/Ben_Cohen_%28businessman%29
Ben Crenshaw	http://en.wikipedia.org/wiki/Ben_Crenshaw
Ben Cross	http://en.wikipedia.org/wiki/Ben_Cross
Ben E. King	http://en.wikipedia.org/wiki/Ben_E._King
Ben Erdreich	http://en.wikipedia.org/wiki/Ben_Erdreich
Ben Folds	http://en.wikipedia.org/wiki/Ben_Folds
Ben Garant	http://en.wikipedia.org/wiki/Ben_Garant
Ben Gazzara	http://en.wikipedia.org/wiki/Ben_Gazzara
Ben Gibbard	http://en.wikipedia.org/wiki/Ben_Gibbard
Ben Harper	http://en.wikipedia.org/wiki/Ben_Harper
Ben Hecht	http://en.wikipedia.org/wiki/Ben_Hecht
Ben Hogan	http://en.wikipedia.org/wiki/Ben_Hogan
Ben Jensen	http://en.wikipedia.org/wiki/Ben_Jensen
Ben Johnson	http://en.wikipedia.org/wiki/Ben_Johnson_%28sprinter%29
Ben Johnson	http://en.wikipedia.org/wiki/Ben_Johnson_%28actor%29
Ben Jones	http://en.wikipedia.org/wiki/Ben_L._Jones
Ben Jonson	http://en.wikipedia.org/wiki/Ben_Jonson
Ben Kingsley	http://en.wikipedia.org/wiki/Ben_Kingsley
Ben Murphy	http://en.wikipedia.org/wiki/Ben_Murphy
Ben Nelson	http://en.wikipedia.org/wiki/Ben_Nelson
Ben Nighthorse Campbell	http://en.wikipedia.org/wiki/Ben_Nighthorse_Campbell
Ben Okri	http://en.wikipedia.org/wiki/Ben_Okri
Ben Pimlott	http://en.wikipedia.org/wiki/Ben_Pimlott
Ben R. Lujan	http://en.wikipedia.org/wiki/Ben_R._Luj%C3%A1n
Ben R. Mottelson	http://en.wikipedia.org/wiki/Ben_R._Mottelson
Ben Roethlisberger	http://en.wikipedia.org/wiki/Ben_Roethlisberger
Ben Savage	http://en.wikipedia.org/wiki/Ben_Savage
Ben Shahn	http://en.wikipedia.org/wiki/Ben_Shahn
Ben Stein	http://en.wikipedia.org/wiki/Ben_Stein
Ben Stiller	http://en.wikipedia.org/wiki/Ben_Stiller
Ben Vereen	http://en.wikipedia.org/wiki/Ben_Vereen
Ben Wallace	http://en.wikipedia.org/wiki/Ben_Wallace
Ben Wallace	http://en.wikipedia.org/wiki/Ben_Wallace_%28UK_politician%29
Ben Wattenberg	http://en.wikipedia.org/wiki/Ben_Wattenberg
Ben Weasel	http://en.wikipedia.org/wiki/Ben_Weasel
Benazir Bhutto	http://en.wikipedia.org/wiki/Benazir_Bhutto
Benedict Arnold	http://en.wikipedia.org/wiki/Benedict_Arnold
Benedict Gummer	http://en.wikipedia.org/wiki/Benedict_Gummer
Benedict XV	http://en.wikipedia.org/wiki/Benedict_XV
Benedict XVI	http://en.wikipedia.org/wiki/Benedict_XVI
Benicio Del Toro	http://en.wikipedia.org/wiki/Benicio_Del_Toro
Benigno Aquino	http://en.wikipedia.org/wiki/Benigno_Aquino_III
Benigno Fitial	http://en.wikipedia.org/wiki/Benigno_Fitial
Benito Mussolini	http://en.wikipedia.org/wiki/Benito_Mussolini
Benjamin A. Gilman	http://en.wikipedia.org/wiki/Benjamin_A._Gilman
Benjamin Apthorp Gould	http://en.wikipedia.org/wiki/Benjamin_Apthorp_Gould
Benjamin Bratt	http://en.wikipedia.org/wiki/Benjamin_Bratt
Benjamin Britten	http://en.wikipedia.org/wiki/Benjamin_Britten
Benjamin Cardozo	http://en.wikipedia.org/wiki/Benjamin_N._Cardozo
Benjamin Count Rumford	http://en.wikipedia.org/wiki/Benjamin_Thompson
Benjamin Disraeli	http://en.wikipedia.org/wiki/Benjamin_Disraeli
Benjamin F. Wade	http://en.wikipedia.org/wiki/Benjamin_F._Wade
Benjamin Franklin	http://en.wikipedia.org/wiki/Benjamin_Franklin
Benjamin Franklin Butler	http://en.wikipedia.org/wiki/Benjamin_Franklin_Butler_%28lawyer%29
Benjamin Harrison	http://en.wikipedia.org/wiki/Benjamin_Harrison
Benjamin Hoadly	http://en.wikipedia.org/wiki/Benjamin_Hoadly
Benjamin Hooks	http://en.wikipedia.org/wiki/Benjamin_Hooks
Benjamin Jowett	http://en.wikipedia.org/wiki/Benjamin_Jowett
Benjamin Kidd	http://en.wikipedia.org/wiki/Benjamin_Kidd
Benjamin L. Cardin	http://en.wikipedia.org/wiki/Benjamin_L._Cardin
Benjamin Latrobe	http://en.wikipedia.org/wiki/Benjamin_Latrobe
Benjamin Lundy	http://en.wikipedia.org/wiki/Benjamin_Lundy
Benjamin McKenzie	http://en.wikipedia.org/wiki/Benjamin_McKenzie
Benjamin Nathaniel Smith	http://en.wikipedia.org/wiki/Benjamin_Nathaniel_Smith
Benjamin Netanyahu	http://en.wikipedia.org/wiki/Benjamin_Netanyahu
Benjamin Orr	http://en.wikipedia.org/wiki/Benjamin_Orr
Benjamin Rush	http://en.wikipedia.org/wiki/Benjamin_Rush
Benjamin Spock	http://en.wikipedia.org/wiki/Benjamin_Spock
Benjamin West	http://en.wikipedia.org/wiki/Benjamin_West
Benji Madden	http://en.wikipedia.org/wiki/Benji_Madden
Bennett Cerf	http://en.wikipedia.org/wiki/Bennett_Cerf
Bennie Thompson	http://en.wikipedia.org/wiki/Bennie_Thompson
Benny Andersen	http://en.wikipedia.org/wiki/Benny_Andersen
Benny Andersson	http://en.wikipedia.org/wiki/Benny_Andersson
Benny Binion	http://en.wikipedia.org/wiki/Benny_Binion
Benny Carter	http://en.wikipedia.org/wiki/Benny_Carter
Benny Goodman	http://en.wikipedia.org/wiki/Benny_Goodman
Benny Hill	http://en.wikipedia.org/wiki/Benny_Hill
Benny Hinn	http://en.wikipedia.org/wiki/Benny_Hinn
Benny Spellman	http://en.wikipedia.org/wiki/Benny_Spellman
Benoit Mandelbrot	http://en.wikipedia.org/wiki/Benoit_Mandelbrot
Benozzo Gozzoli	http://en.wikipedia.org/wiki/Benozzo_Gozzoli
Benvenuto Cellini	http://en.wikipedia.org/wiki/Benvenuto_Cellini
Berengar of Tours	http://en.wikipedia.org/wiki/Berengar_of_Tours
Berke Breathed	http://en.wikipedia.org/wiki/Berke_Breathed
Berkley Bedell	http://en.wikipedia.org/wiki/Berkley_Bedell
Bern Nadette Stanis	http://en.wikipedia.org/wiki/Bern_Nadette_Stanis
Bernadette Devlin	http://en.wikipedia.org/wiki/Bernadette_Devlin_McAliskey
Bernadette Peters	http://en.wikipedia.org/wiki/Bernadette_Peters
Bernard Addison	http://en.wikipedia.org/wiki/Bernard_Addison
Bernard Arnault	http://en.wikipedia.org/wiki/Bernard_Arnault
Bernard Cornwell	http://en.wikipedia.org/wiki/Bernard_Cornwell
Bernard de Mandeville	http://en.wikipedia.org/wiki/Bernard_de_Mandeville
Bernard Ebbers	http://en.wikipedia.org/wiki/Bernard_Ebbers
Bernard Edwards	http://en.wikipedia.org/wiki/Bernard_Edwards
Bernard Goldberg	http://en.wikipedia.org/wiki/Bernard_Goldberg
Bernard Herrmann	http://en.wikipedia.org/wiki/Bernard_Herrmann
Bernard Hill	http://en.wikipedia.org/wiki/Bernard_Hill
Bernard J. Dwyer	http://en.wikipedia.org/wiki/Bernard_J._Dwyer
Bernard Jenkin	http://en.wikipedia.org/wiki/Bernard_Jenkin
Bernard Kalb	http://en.wikipedia.org/wiki/Bernard_Kalb
Bernard Kerik	http://en.wikipedia.org/wiki/Bernard_Kerik
Bernard Law	http://en.wikipedia.org/wiki/Bernard_Law
Bernard le Bovier de Fontenelle	http://en.wikipedia.org/wiki/Bernard_le_Bovier_de_Fontenelle
Bernard Lee	http://en.wikipedia.org/wiki/Bernard_Lee
Bernard Lintot	http://en.wikipedia.org/wiki/Bernard_Lintot
Bernard M. Baruch	http://en.wikipedia.org/wiki/Bernard_M._Baruch
Bernard Makuza	http://en.wikipedia.org/wiki/Bernard_Makuza
Bernard Malamud	http://en.wikipedia.org/wiki/Bernard_Malamud
Bernard Montgomery	http://en.wikipedia.org/wiki/Bernard_Montgomery
Bernard Shaw	http://en.wikipedia.org/wiki/Bernard_Shaw_%28journalist%29
Bernard Sumner	http://en.wikipedia.org/wiki/Bernard_Sumner
Bernard Trainor	http://en.wikipedia.org/wiki/Bernard_Trainor
Bernard van Orley	http://en.wikipedia.org/wiki/Bernard_van_Orley
Bernard-Henri L�vy	http://en.wikipedia.org/wiki/Bernard-Henri_L%C3%A9vy
Bernardim Ribeiro	http://en.wikipedia.org/wiki/Bernardim_Ribeiro
Bernardino Luini	http://en.wikipedia.org/wiki/Bernardino_Luini
Bernardino Telesio	http://en.wikipedia.org/wiki/Bernardino_Telesio
Bernardo Bertolucci	http://en.wikipedia.org/wiki/Bernardo_Bertolucci
Bernardo O'Higgins	http://en.wikipedia.org/wiki/Bernardo_O%27Higgins
Bernhard Goetz	http://en.wikipedia.org/wiki/Bernhard_Goetz
Bernhard Riemann	http://en.wikipedia.org/wiki/Bernhard_Riemann
Bernhard von Bulow	http://en.wikipedia.org/wiki/Bernhard_von_Bulow
Bernie Allen	http://en.wikipedia.org/wiki/Bernie_Allen
Bernie Casey	http://en.wikipedia.org/wiki/Bernie_Casey
Bernie Kopell	http://en.wikipedia.org/wiki/Bernie_Kopell
Bernie Krause	http://en.wikipedia.org/wiki/Bernie_Krause
Bernie Mac	http://en.wikipedia.org/wiki/Bernie_Mac
Bernie Sanders	http://en.wikipedia.org/wiki/Bernie_Sanders
Bernie Taupin	http://en.wikipedia.org/wiki/Bernie_Taupin
Bernie Ward	http://en.wikipedia.org/wiki/Bernie_Ward
Bernie Worrell	http://en.wikipedia.org/wiki/Bernie_Worrell
Berry Gordy	http://en.wikipedia.org/wiki/Berry_Gordy
Bert Campaneris	http://en.wikipedia.org/wiki/Bert_Campaneris
Bert Convy	http://en.wikipedia.org/wiki/Bert_Convy
Bert I. Gordon	http://en.wikipedia.org/wiki/Bert_I._Gordon
Bert Lahr	http://en.wikipedia.org/wiki/Bert_Lahr
Bert McCracken	http://en.wikipedia.org/wiki/Bert_McCracken
Bert Parks	http://en.wikipedia.org/wiki/Bert_Parks
Bertha von Suttner	http://en.wikipedia.org/wiki/Bertha_von_Suttner
Berthe Morisot	http://en.wikipedia.org/wiki/Berthe_Morisot
Bertie Ahern	http://en.wikipedia.org/wiki/Bertie_Ahern
Bertie Forbes	http://en.wikipedia.org/wiki/Bertie_Forbes
Bertil Ohlin	http://en.wikipedia.org/wiki/Bertil_Ohlin
Bertolt Brecht	http://en.wikipedia.org/wiki/Bertolt_Brecht
Bertram N. Brockhouse	http://en.wikipedia.org/wiki/Bertram_N._Brockhouse
Bertrand Cantat	http://en.wikipedia.org/wiki/Bertrand_Cantat
Bertrand H. Snell	http://en.wikipedia.org/wiki/Bertrand_H._Snell
Bertrand R. Brinley	http://en.wikipedia.org/wiki/Bertrand_R._Brinley
Bertrand Russell	http://en.wikipedia.org/wiki/Bertrand_Russell
Beryl Anthony, Jr.	http://en.wikipedia.org/wiki/Beryl_Anthony,_Jr.
Beryl Bainbridge	http://en.wikipedia.org/wiki/Beryl_Bainbridge
Bess Armstrong	http://en.wikipedia.org/wiki/Bess_Armstrong
Bess Myerson	http://en.wikipedia.org/wiki/Bess_Myerson
Bess Truman	http://en.wikipedia.org/wiki/Bess_Truman
Bessie Head	http://en.wikipedia.org/wiki/Bessie_Head
Bessie Love	http://en.wikipedia.org/wiki/Bessie_Love
Bessie Potter Vonnoh	http://en.wikipedia.org/wiki/Bessie_Potter_Vonnoh
Bessie Smith	http://en.wikipedia.org/wiki/Bessie_Smith
Beth Allen	http://en.wikipedia.org/wiki/Beth_Allen
Beth Gibbons	http://en.wikipedia.org/wiki/Beth_Gibbons
Beth Henley	http://en.wikipedia.org/wiki/Beth_Henley
Beth Orton	http://en.wikipedia.org/wiki/Beth_Orton
Beth Ostrosky	http://en.wikipedia.org/wiki/Beth_Ostrosky
Bethany Joy Lenz	http://en.wikipedia.org/wiki/Bethany_Joy_Lenz
Betsy Markey	http://en.wikipedia.org/wiki/Betsy_Markey
Betsy Palmer	http://en.wikipedia.org/wiki/Betsy_Palmer
Betsy Ross	http://en.wikipedia.org/wiki/Betsy_Ross
Bette Davis	http://en.wikipedia.org/wiki/Bette_Davis
Bette Midler	http://en.wikipedia.org/wiki/Bette_Midler
Bettie Page	http://en.wikipedia.org/wiki/Bettie_Page
Bettino Craxi	http://en.wikipedia.org/wiki/Bettino_Craxi
Betty Buckley	http://en.wikipedia.org/wiki/Betty_Buckley
Betty Dodson	http://en.wikipedia.org/wiki/Betty_Dodson
Betty Ford	http://en.wikipedia.org/wiki/Betty_Ford
Betty Friedan	http://en.wikipedia.org/wiki/Betty_Friedan
Betty Grable	http://en.wikipedia.org/wiki/Betty_Grable
Betty Hill	http://en.wikipedia.org/wiki/Betty_Hill
Betty Hutton	http://en.wikipedia.org/wiki/Betty_Hutton
Betty McCollum	http://en.wikipedia.org/wiki/Betty_McCollum
Betty Shabazz	http://en.wikipedia.org/wiki/Betty_Shabazz
Betty Smith	http://en.wikipedia.org/wiki/Betty_Smith
Betty Sutton	http://en.wikipedia.org/wiki/Betty_Sutton
Betty Thomas	http://en.wikipedia.org/wiki/Betty_Thomas
Betty White	http://en.wikipedia.org/wiki/Betty_White
Betty Williams	http://en.wikipedia.org/wiki/Betty_Williams_%28Nobel_laureate%29
Bev Bevan	http://en.wikipedia.org/wiki/Bev_Bevan
Beverley Mitchell	http://en.wikipedia.org/wiki/Beverley_Mitchell
Beverly B. Byron	http://en.wikipedia.org/wiki/Beverly_B._Byron
Beverly Cleary	http://en.wikipedia.org/wiki/Beverly_Cleary
Beverly D'Angelo	http://en.wikipedia.org/wiki/Beverly_D%27Angelo
Beverly LaHaye	http://en.wikipedia.org/wiki/Beverly_LaHaye
Beverly Sills	http://en.wikipedia.org/wiki/Beverly_Sills
Beyonce Knowles	http://en.wikipedia.org/wiki/Beyonce_Knowles
Bhagwan Shree Rajneesh	http://en.wikipedia.org/wiki/Bhagwan_Shree_Rajneesh
Bharati Mukherjee	http://en.wikipedia.org/wiki/Bharati_Mukherjee
Bharrat Jagdeo	http://en.wikipedia.org/wiki/Bharrat_Jagdeo
Bhumibol Adulyadej	http://en.wikipedia.org/wiki/Bhumibol_Adulyadej
Bianca Jagger	http://en.wikipedia.org/wiki/Bianca_Jagger
Bibbe Hansen	http://en.wikipedia.org/wiki/Bibbe_Hansen
Bibi Besch	http://en.wikipedia.org/wiki/Bibi_Besch
Big Boi	http://en.wikipedia.org/wiki/Big_Boi
Big Daddy Kane	http://en.wikipedia.org/wiki/Big_Daddy_Kane
Big Joe Turner	http://en.wikipedia.org/wiki/Big_Joe_Turner
Big Pun	http://en.wikipedia.org/wiki/Big_Pun
Bijou Phillips	http://en.wikipedia.org/wiki/Bijou_Phillips
Bil Keane	http://en.wikipedia.org/wiki/Bil_Keane
Bill Archer	http://en.wikipedia.org/wiki/William_Reynolds_Archer,_Jr.
Bill Arp	http://en.wikipedia.org/wiki/Bill_Arp
Bill Ballance	http://en.wikipedia.org/wiki/Bill_Ballance
Bill Bass	http://en.wikipedia.org/wiki/Bill_Bass
Bill Bellamy	http://en.wikipedia.org/wiki/Bill_Bellamy
Bill Bixby	http://en.wikipedia.org/wiki/Bill_Bixby
Bill Blass	http://en.wikipedia.org/wiki/Bill_Blass
Bill Boner	http://en.wikipedia.org/wiki/Bill_Boner
Bill Bradley	http://en.wikipedia.org/wiki/Bill_Bradley
Bill Bruford	http://en.wikipedia.org/wiki/Bill_Bruford
Bill Buckner	http://en.wikipedia.org/wiki/Bill_Buckner
Bill Budge	http://en.wikipedia.org/wiki/Bill_Budge
Bill Callahan	http://en.wikipedia.org/wiki/Bill_Callahan_%28musician%29
Bill Campbell	http://en.wikipedia.org/wiki/Bill_Campbell_%28mayor%29
Bill Cassidy	http://en.wikipedia.org/wiki/Bill_Cassidy
Bill Clinton	http://en.wikipedia.org/wiki/Bill_Clinton
Bill Cobey	http://en.wikipedia.org/wiki/Bill_Cobey
Bill Condon	http://en.wikipedia.org/wiki/Bill_Condon
Bill Cosby	http://en.wikipedia.org/wiki/Bill_Cosby
Bill Cullen	http://en.wikipedia.org/wiki/Bill_Cullen
Bill Daily	http://en.wikipedia.org/wiki/Bill_Daily
Bill Delahunt	http://en.wikipedia.org/wiki/Bill_Delahunt
Bill Dickey	http://en.wikipedia.org/wiki/Bill_Dickey
Bill Dickinson	http://en.wikipedia.org/wiki/William_Louis_Dickinson
Bill Donaldson	http://en.wikipedia.org/wiki/Bill_Donaldson
Bill Emerson	http://en.wikipedia.org/wiki/Bill_Emerson
Bill Esterson	http://en.wikipedia.org/wiki/Bill_Esterson
Bill Foster	http://en.wikipedia.org/wiki/Bill_Foster_%28Illinois_politician%29
Bill France, Jr.	http://en.wikipedia.org/wiki/Bill_France,_Jr.
Bill Frenzel	http://en.wikipedia.org/wiki/Bill_Frenzel
Bill Frisell	http://en.wikipedia.org/wiki/Bill_Frisell
Bill Frist	http://en.wikipedia.org/wiki/Bill_Frist
Bill Gates	http://en.wikipedia.org/wiki/Bill_Gates
Bill Geist	http://en.wikipedia.org/wiki/Bill_Geist
Bill Gertz	http://en.wikipedia.org/wiki/Bill_Gertz
Bill Goldberg	http://en.wikipedia.org/wiki/Bill_Goldberg
Bill Graham	http://en.wikipedia.org/wiki/Bill_Graham
Bill Griffith	http://en.wikipedia.org/wiki/Bill_Griffith
Bill Haley	http://en.wikipedia.org/wiki/Bill_Haley
Bill Hefner	http://en.wikipedia.org/wiki/Bill_Hefner
Bill Hemmer	http://en.wikipedia.org/wiki/Bill_Hemmer
Bill Hendon	http://en.wikipedia.org/wiki/Bill_Hendon
Bill Hicks	http://en.wikipedia.org/wiki/Bill_Hicks
Bill Janklow	http://en.wikipedia.org/wiki/Bill_Janklow
Bill Joy	http://en.wikipedia.org/wiki/Bill_Joy
Bill Justis	http://en.wikipedia.org/wiki/Bill_Justis
Bill Keller	http://en.wikipedia.org/wiki/Bill_Keller
Bill Kreutzman	http://en.wikipedia.org/wiki/Bill_Kreutzman
Bill Kristol	http://en.wikipedia.org/wiki/Bill_Kristol
Bill Kurtis	http://en.wikipedia.org/wiki/Bill_Kurtis
Bill Laimbeer	http://en.wikipedia.org/wiki/Bill_Laimbeer
Bill Laswell	http://en.wikipedia.org/wiki/Bill_Laswell
Bill Lipinski	http://en.wikipedia.org/wiki/Bill_Lipinski
Bill Lowery	http://en.wikipedia.org/wiki/Bill_Lowery
Bill Luther	http://en.wikipedia.org/wiki/Bill_Luther
Bill Macy	http://en.wikipedia.org/wiki/Bill_Macy
Bill Maher	http://en.wikipedia.org/wiki/Bill_Maher
Bill Mazeroski	http://en.wikipedia.org/wiki/Bill_Mazeroski
Bill McCollum	http://en.wikipedia.org/wiki/Bill_McCollum
Bill Melendez	http://en.wikipedia.org/wiki/Bill_Melendez
Bill Morrow	http://en.wikipedia.org/wiki/Bill_Morrow_%28California_politician%29
Bill Moyers	http://en.wikipedia.org/wiki/Bill_Moyers
Bill Mumy	http://en.wikipedia.org/wiki/Bill_Mumy
Bill Murray	http://en.wikipedia.org/wiki/Bill_Murray
Bill Nelson	http://en.wikipedia.org/wiki/Bill_Nelson
Bill Nichols	http://en.wikipedia.org/wiki/William_Flynt_Nichols
Bill Nighy	http://en.wikipedia.org/wiki/Bill_Nighy
Bill Nye	http://en.wikipedia.org/wiki/Bill_Nye
Bill Nye	http://en.wikipedia.org/wiki/Edgar_Wilson_Nye
Bill O'Reilly	http://en.wikipedia.org/wiki/Bill_O%27Reilly_%28political_commentator%29
Bill Owen	http://en.wikipedia.org/wiki/Bill_Owen_%28actor%29
Bill Owens	http://en.wikipedia.org/wiki/Bill_Owens_%28Colorado_politician%29
Bill Owens	http://en.wikipedia.org/wiki/Bill_Owens_%28congressman%29
Bill Parcells	http://en.wikipedia.org/wiki/Bill_Parcells
Bill Pascrell	http://en.wikipedia.org/wiki/Bill_Pascrell
Bill Paxton	http://en.wikipedia.org/wiki/Bill_Paxton
Bill Pearl	http://en.wikipedia.org/wiki/Bill_Pearl
Bill Posey	http://en.wikipedia.org/wiki/Bill_Posey
Bill Pullman	http://en.wikipedia.org/wiki/Bill_Pullman
Bill Richardson	http://en.wikipedia.org/wiki/Bill_Richardson
Bill Romanowski	http://en.wikipedia.org/wiki/Bill_Romanowski
Bill Russell	http://en.wikipedia.org/wiki/Bill_Russell
Bill Saluga	http://en.wikipedia.org/wiki/Bill_Saluga
Bill Schneider	http://en.wikipedia.org/wiki/Bill_Schneider_%28journalist%29
Bill Schuette	http://en.wikipedia.org/wiki/Bill_Schuette
Bill Scott	http://en.wikipedia.org/wiki/Bill_Scott_%28voice_actor%29
Bill Shankly	http://en.wikipedia.org/wiki/Bill_Shankly
Bill Sharman	http://en.wikipedia.org/wiki/Bill_Sharman
Bill Shuster	http://en.wikipedia.org/wiki/Bill_Shuster
Bill Sienkiewicz	http://en.wikipedia.org/wiki/Bill_Sienkiewicz
Bill Thomas	http://en.wikipedia.org/wiki/Bill_Thomas
Bill Veeck	http://en.wikipedia.org/wiki/Bill_Veeck
Bill Walton	http://en.wikipedia.org/wiki/Bill_Walton
Bill Ward	http://en.wikipedia.org/wiki/Bill_Ward_%28musician%29
Bill Watterson	http://en.wikipedia.org/wiki/Bill_Watterson
Bill Weld	http://en.wikipedia.org/wiki/Bill_Weld
Bill Wiggin	http://en.wikipedia.org/wiki/Bill_Wiggin
Bill Williams	http://en.wikipedia.org/wiki/Bill_Williams_%28actor%29
Bill Wyman	http://en.wikipedia.org/wiki/Bill_Wyman
Bill Young	http://en.wikipedia.org/wiki/Bill_Young
Bille August	http://en.wikipedia.org/wiki/Bille_August
Bille Jean King	http://en.wikipedia.org/wiki/Billie_Jean_King
Billie Burke	http://en.wikipedia.org/wiki/Billie_Burke
Billie Holiday	http://en.wikipedia.org/wiki/Billie_Holiday
Billie Joe Armstrong	http://en.wikipedia.org/wiki/Billie_Joe_Armstrong
Billie Piper	http://en.wikipedia.org/wiki/Billie_Piper
Billy Barty	http://en.wikipedia.org/wiki/Billy_Barty
Billy Bean	http://en.wikipedia.org/wiki/Billy_Bean
Billy Beane	http://en.wikipedia.org/wiki/Billy_Beane
Billy Blanks	http://en.wikipedia.org/wiki/Billy_Blanks
Billy Bob Thornton	http://en.wikipedia.org/wiki/Billy_Bob_Thornton
Billy Boyd	http://en.wikipedia.org/wiki/Billy_Boyd_%28actor%29
Billy Bragg	http://en.wikipedia.org/wiki/Billy_Bragg
Billy Bush	http://en.wikipedia.org/wiki/Billy_Bush
Billy Campbell	http://en.wikipedia.org/wiki/Billy_Campbell
Billy Carter	http://en.wikipedia.org/wiki/Billy_Carter
Billy Connolly	http://en.wikipedia.org/wiki/Billy_Connolly
Billy Corgan	http://en.wikipedia.org/wiki/Billy_Corgan
Billy Crudup	http://en.wikipedia.org/wiki/Billy_Crudup
Billy Crystal	http://en.wikipedia.org/wiki/Billy_Crystal
Billy Dee Williams	http://en.wikipedia.org/wiki/Billy_Dee_Williams
Billy Drago	http://en.wikipedia.org/wiki/Billy_Drago
Billy Eckstine	http://en.wikipedia.org/wiki/Billy_Eckstine
Billy Fury	http://en.wikipedia.org/wiki/Billy_Fury
Billy Graham	http://en.wikipedia.org/wiki/Billy_Graham
Billy Gray	http://en.wikipedia.org/wiki/Billy_Gray
Billy Higgins	http://en.wikipedia.org/wiki/Billy_Higgins
Billy Howerdel	http://en.wikipedia.org/wiki/Billy_Howerdel
Billy Idol	http://en.wikipedia.org/wiki/Billy_Idol
Billy Joel	http://en.wikipedia.org/wiki/Billy_Joel
Billy Kl�ver	http://en.wikipedia.org/wiki/Billy_Kl%C3%Bcver
Billy Martin	http://en.wikipedia.org/wiki/Billy_Martin_%28guitarist%29
Billy Martin	http://en.wikipedia.org/wiki/Billy_Martin
Billy Mays 	http://en.wikipedia.org/wiki/Billy_mays
Billy Morrison	http://en.wikipedia.org/wiki/Billy_Morrison
Billy Murray	http://en.wikipedia.org/wiki/Billy_Murray_%28singer%29
Billy Ocean	http://en.wikipedia.org/wiki/Billy_Ocean
Billy Powell	http://en.wikipedia.org/wiki/Billy_Powell
Billy Preston	http://en.wikipedia.org/wiki/Billy_Preston
Billy Ray Cyrus	http://en.wikipedia.org/wiki/Billy_Ray_Cyrus
Billy Sheehan	http://en.wikipedia.org/wiki/Billy_Sheehan
Billy Sherwood	http://en.wikipedia.org/wiki/Billy_Sherwood
Billy Sims	http://en.wikipedia.org/wiki/Billy_Sims
Billy Squier	http://en.wikipedia.org/wiki/Billy_Squier
Billy Tauzin	http://en.wikipedia.org/wiki/Billy_Tauzin
Billy the Kid	http://en.wikipedia.org/wiki/Billy_the_Kid
Billy Thorpe	http://en.wikipedia.org/wiki/Billy_Thorpe
Billy West	http://en.wikipedia.org/wiki/Billy_West
Billy Wilder	http://en.wikipedia.org/wiki/Billy_Wilder
Billy Williams	http://en.wikipedia.org/wiki/Billy_Williams_%28baseball%29
Billy Zane	http://en.wikipedia.org/wiki/Billy_Zane
Bing Crosby	http://en.wikipedia.org/wiki/Bing_Crosby
Bingu wa Mutharika	http://en.wikipedia.org/wiki/Bingu_wa_Mutharika
Birch Bayh	http://en.wikipedia.org/wiki/Birch_Bayh
Bird McIntyre	http://en.wikipedia.org/wiki/Bird_McIntyre
Birdman of Alcatraz	http://en.wikipedia.org/wiki/Birdman_of_Alcatraz
Birgit Nilsson	http://en.wikipedia.org/wiki/Birgit_Nilsson
Birut Galdikas	http://en.wikipedia.org/wiki/Birut%C3%A9_Galdikas
Bix Beiderbecke	http://en.wikipedia.org/wiki/Bix_Beiderbecke
Biz Markie	http://en.wikipedia.org/wiki/Biz_Markie
Bizzy Bone	http://en.wikipedia.org/wiki/Bizzy_Bone
Bjarne Stroustrup	http://en.wikipedia.org/wiki/Bjarne_Stroustrup
Bjorn Borg	http://en.wikipedia.org/wiki/Bjorn_Borg
Bj�rn Lomborg	http://en.wikipedia.org/wiki/Bj%C3%B8rn_Lomborg
Bj�rn Ulvaeus	http://en.wikipedia.org/wiki/Bj%C3%B6rn_Ulvaeus
Blackie Lawless	http://en.wikipedia.org/wiki/Blackie_Lawless
Blag Dahlia	http://en.wikipedia.org/wiki/Blag_Dahlia
Blaine Luetkemeyer	http://en.wikipedia.org/wiki/Blaine_Luetkemeyer
Blair Brown	http://en.wikipedia.org/wiki/Blair_Brown
Blair Underwood	http://en.wikipedia.org/wiki/Blair_Underwood
Blaise Compaor�	http://en.wikipedia.org/wiki/Blaise_Compaor%c3%a9
Blaise Pascal	http://en.wikipedia.org/wiki/Blaise_Pascal
Blake Edwards	http://en.wikipedia.org/wiki/Blake_Edwards
Blake Lively	http://en.wikipedia.org/wiki/Blake_Lively
Blanche Lincoln	http://en.wikipedia.org/wiki/Blanche_Lincoln
Blaze Starr	http://en.wikipedia.org/wiki/Blaze_Starr
Blessed John XXIII	http://en.wikipedia.org/wiki/Blessed_John_XXIII
Blind Harry	http://en.wikipedia.org/wiki/Blind_Harry
Blixa Bargeld	http://en.wikipedia.org/wiki/Blixa_Bargeld
Blythe Danner	http://en.wikipedia.org/wiki/Blythe_Danner
Bo Bice	http://en.wikipedia.org/wiki/Bo_Bice
Bo Derek	http://en.wikipedia.org/wiki/Bo_Derek
Bo Diddley	http://en.wikipedia.org/wiki/Bo_Diddley
Bo Dietl	http://en.wikipedia.org/wiki/Bo_Dietl
Bo Gritz	http://en.wikipedia.org/wiki/Bo_Gritz
Bo Hi Pak	http://en.wikipedia.org/wiki/Bo_Hi_Pak
Bo Jackson	http://en.wikipedia.org/wiki/Bo_Jackson
Bob Abernethy	http://en.wikipedia.org/wiki/Bob_Abernethy
Bob Adrian	http://en.wikipedia.org/wiki/Bob_Adrian
Bob Ainsworth	http://en.wikipedia.org/wiki/Bob_Ainsworth
Bob Allen	http://en.wikipedia.org/wiki/Bob_Allen
Bob Balaban	http://en.wikipedia.org/wiki/Bob_Balaban
Bob Barker	http://en.wikipedia.org/wiki/Bob_Barker
Bob Barr	http://en.wikipedia.org/wiki/Bob_Barr
Bob Beauprez	http://en.wikipedia.org/wiki/Bob_Beauprez
Bob Blackman	http://en.wikipedia.org/wiki/Robert_Blackman
Bob Brinker	http://en.wikipedia.org/wiki/Bob_Brinker
Bob Bryar	http://en.wikipedia.org/wiki/Bob_Bryar
Bob Burns	http://en.wikipedia.org/wiki/Bob_Burns_%28politician%29
Bob Carr	http://en.wikipedia.org/wiki/Bob_Carr
Bob Clement	http://en.wikipedia.org/wiki/Bob_Clement
Bob Corker	http://en.wikipedia.org/wiki/Bob_Corker
Bob Costas	http://en.wikipedia.org/wiki/Bob_Costas
Bob Cousy	http://en.wikipedia.org/wiki/Bob_Cousy
Bob Crane	http://en.wikipedia.org/wiki/Bob_Crane
Bob Cummings	http://en.wikipedia.org/wiki/Bob_Cummings
Bob Denver	http://en.wikipedia.org/wiki/Bob_Denver
Bob Dole	http://en.wikipedia.org/wiki/Bob_Dole
Bob Dornan	http://en.wikipedia.org/wiki/Bob_Dornan
Bob Dylan	http://en.wikipedia.org/wiki/Bob_Dylan
Bob Edgar	http://en.wikipedia.org/wiki/Bob_Edgar
Bob Edwards	http://en.wikipedia.org/wiki/Bob_Edwards
Bob Elliott	http://en.wikipedia.org/wiki/Bob_Elliott_%28basketball%29
Bob Etheridge	http://en.wikipedia.org/wiki/Bob_Etheridge
Bob Eubanks	http://en.wikipedia.org/wiki/Bob_Eubanks
Bob Feller	http://en.wikipedia.org/wiki/Bob_Feller
Bob Filner	http://en.wikipedia.org/wiki/Bob_Filner
Bob Fosse	http://en.wikipedia.org/wiki/Bob_Fosse
Bob Franks	http://en.wikipedia.org/wiki/Bob_Franks
Bob Frankston	http://en.wikipedia.org/wiki/Bob_Frankston
Bob Geldof	http://en.wikipedia.org/wiki/Bob_Geldof
Bob Gibson	http://en.wikipedia.org/wiki/Bob_Gibson
Bob Goldthwait	http://en.wikipedia.org/wiki/Bob_Goldthwait
Bob Goodlatte	http://en.wikipedia.org/wiki/Bob_Goodlatte
Bob Graham	http://en.wikipedia.org/wiki/Bob_Graham
Bob Grant	http://en.wikipedia.org/wiki/Bob_Grant_%28radio%29
Bob Griese	http://en.wikipedia.org/wiki/Bob_Griese
Bob Guccione	http://en.wikipedia.org/wiki/Bob_Guccione
Bob Guccione, Jr.	http://en.wikipedia.org/wiki/Bob_Guccione,_Jr.
Bob Holden	http://en.wikipedia.org/wiki/Bob_Holden
Bob Hope	http://en.wikipedia.org/wiki/Bob_Hope
Bob Hoskins	http://en.wikipedia.org/wiki/Bob_Hoskins
Bob Inglis	http://en.wikipedia.org/wiki/Bob_Inglis
Bob Irwin	http://en.wikipedia.org/wiki/Bob_Irwin
Bob Kane	http://en.wikipedia.org/wiki/Bob_Kane
Bob Kasten	http://en.wikipedia.org/wiki/Bob_Kasten
Bob Kaufman	http://en.wikipedia.org/wiki/Bob_Kaufman
Bob Kerrey	http://en.wikipedia.org/wiki/Bob_Kerrey
Bob Latta	http://en.wikipedia.org/wiki/Bob_Latta
Bob Livingston	http://en.wikipedia.org/wiki/Bob_Livingston
Bob Mackie	http://en.wikipedia.org/wiki/Bob_Mackie
Bob Marley	http://en.wikipedia.org/wiki/Bob_Marley
Bob Mathias	http://en.wikipedia.org/wiki/Bob_Mathias
Bob McAdoo	http://en.wikipedia.org/wiki/Bob_McAdoo
Bob Menendez	http://en.wikipedia.org/wiki/Bob_Menendez
Bob Metcalfe	http://en.wikipedia.org/wiki/Bob_Metcalfe
Bob Miller	http://en.wikipedia.org/wiki/Rob_Miller_%28South_Carolina_politician%29
Bob Mould	http://en.wikipedia.org/wiki/Bob_Mould
Bob Neill	http://en.wikipedia.org/wiki/Bob_Neill
Bob Newhart	http://en.wikipedia.org/wiki/Bob_Newhart
Bob Ney	http://en.wikipedia.org/wiki/Bob_Ney
Bob Odenkirk	http://en.wikipedia.org/wiki/Bob_Odenkirk
Bob Packwood	http://en.wikipedia.org/wiki/Bob_Packwood
Bob Paisley	http://en.wikipedia.org/wiki/Bob_Paisley
Bob Pettit	http://en.wikipedia.org/wiki/Bob_Pettit
Bob Probert	http://en.wikipedia.org/wiki/Bob_Probert
Bob Rafelson	http://en.wikipedia.org/wiki/Bob_Rafelson
Bob Riley	http://en.wikipedia.org/wiki/Bob_Riley
Bob Ross	http://en.wikipedia.org/wiki/Bob_Ross
Bob Russell	http://en.wikipedia.org/wiki/Bob_Russell_%28politician%29
Bob Saget	http://en.wikipedia.org/wiki/Bob_Saget
Bob Schaffer	http://en.wikipedia.org/wiki/Bob_Schaffer
Bob Schieffer	http://en.wikipedia.org/wiki/Bob_Schieffer
Bob Seger	http://en.wikipedia.org/wiki/Bob_Seger
Bob Shaw	http://en.wikipedia.org/wiki/Bob_Shaw
Bob Simon	http://en.wikipedia.org/wiki/Bob_Simon
Bob Smith	http://en.wikipedia.org/wiki/Bob_Smith_%28New_Jersey_State_Senator%29
Bob Somerby	http://en.wikipedia.org/wiki/Bob_Somerby
Bob Stanley	http://en.wikipedia.org/wiki/Bob_Stanley
Bob Stewart	http://en.wikipedia.org/wiki/Bob_Stewart_(British_Army_officer)
Bob Stump	http://en.wikipedia.org/wiki/Bob_Stump
Bob Taft	http://en.wikipedia.org/wiki/Bob_Taft
Bob Tisch	http://en.wikipedia.org/wiki/Bob_Tisch
Bob Traxler	http://en.wikipedia.org/wiki/Bob_Traxler
Bob Uecker	http://en.wikipedia.org/wiki/Bob_Uecker
Bob Vila	http://en.wikipedia.org/wiki/Bob_Vila
Bob Weir	http://en.wikipedia.org/wiki/Bob_Weir
Bob West	http://en.wikipedia.org/wiki/Bob_West
Bob Whittaker	http://en.wikipedia.org/wiki/Bob_Whittaker
Bob Wise	http://en.wikipedia.org/wiki/Bob_Wise
Bob Woodruff	http://en.wikipedia.org/wiki/Bob_Woodruff
Bob Woodward	http://en.wikipedia.org/wiki/Bob_Woodward
Bobbi Fiedler	http://en.wikipedia.org/wiki/Bobbi_Fiedler
Bobbie Ann Mason	http://en.wikipedia.org/wiki/Bobbie_Ann_Mason
Bobbie Gentry	http://en.wikipedia.org/wiki/Bobbie_Gentry
Bobby "The Brain" Heenan	http://en.wikipedia.org/wiki/Bobby_%22The_Brain%22_Heenan
Bobby Allen	http://en.wikipedia.org/wiki/Bobby_Allen
Bobby Bland	http://en.wikipedia.org/wiki/Bobby_Bland
Bobby Bonilla	http://en.wikipedia.org/wiki/Bobby_Bonilla
Bobby Bowden	http://en.wikipedia.org/wiki/Bobby_Bowden
Bobby Bright	http://en.wikipedia.org/wiki/Bobby_Bright
Bobby Brown	http://en.wikipedia.org/wiki/Bobby_Brown
Bobby Cannavale	http://en.wikipedia.org/wiki/Bobby_Cannavale
Bobby Charlton	http://en.wikipedia.org/wiki/Bobby_Charlton
Bobby Darin	http://en.wikipedia.org/wiki/Bobby_Darin
Bobby Day	http://en.wikipedia.org/wiki/Bobby_Day
Bobby Driscoll	http://en.wikipedia.org/wiki/Bobby_Driscoll
Bobby Edner	http://en.wikipedia.org/wiki/Bobby_Edner
Bobby Farrelly	http://en.wikipedia.org/wiki/Bobby_Farrelly
Bobby Fischer	http://en.wikipedia.org/wiki/Bobby_Fischer
Bobby Flay	http://en.wikipedia.org/wiki/Bobby_Flay
Bobby Gillespie	http://en.wikipedia.org/wiki/Bobby_Gillespie
Bobby Hull	http://en.wikipedia.org/wiki/Bobby_Hull
Bobby Jindal	http://en.wikipedia.org/wiki/Bobby_Jindal
Bobby Jones	http://en.wikipedia.org/wiki/Bobby_Jones_(golfer)
Bobby Kimball	http://en.wikipedia.org/wiki/Bobby_Kimball
Bobby Knight	http://en.wikipedia.org/wiki/Bobby_Knight
Bobby McFerrin	http://en.wikipedia.org/wiki/Bobby_McFerrin
Bobby Moore	http://en.wikipedia.org/wiki/Bobby_Moore
Bobby Orr	http://en.wikipedia.org/wiki/Bobby_Orr
Bobby Rahal	http://en.wikipedia.org/wiki/Bobby_Rahal
Bobby Ray Inman	http://en.wikipedia.org/wiki/Bobby_Ray_Inman
Bobby Rush	http://en.wikipedia.org/wiki/Bobby_Rush
Bobby Sands	http://en.wikipedia.org/wiki/Bobby_Sands
Bobby Scott	http://en.wikipedia.org/wiki/Robert_C._Scott
Bobby Seale	http://en.wikipedia.org/wiki/Bobby_Seale
Bobby Sherman	http://en.wikipedia.org/wiki/Bobby_Sherman
Bobby Short	http://en.wikipedia.org/wiki/Bobby_Short
Bobby Shriver	http://en.wikipedia.org/wiki/Bobby_Shriver
Bobby Thomson	http://en.wikipedia.org/wiki/Bobby_Thomson
Bobby Trendy	http://en.wikipedia.org/wiki/Bobby_Trendy
Bobby Unser	http://en.wikipedia.org/wiki/Bobby_Unser
Bobby Valentino	http://en.wikipedia.org/wiki/Bobby_Valentino
Bobby Vinton	http://en.wikipedia.org/wiki/Bobby_Vinton
Bobby Womack	http://en.wikipedia.org/wiki/Bobby_Womack
Bobcat Goldthwait	http://en.wikipedia.org/wiki/Bobcat_Goldthwait
Bodhi Elfman	http://en.wikipedia.org/wiki/Bodhi_Elfman
Bogdan Raczynski	http://en.wikipedia.org/wiki/Bogdan_Raczynski
Bohumil Hrabal	http://en.wikipedia.org/wiki/Bohumil_Hrabal
Bojan Kostreš	http://en.wikipedia.org/wiki/Bojan_Kostre%C5%A1
Bojan Pajtic	http://en.wikipedia.org/wiki/Bojan_Pajtic
Bon Scott	http://en.wikipedia.org/wiki/Bon_Scott
Bonaventure des P�riers	http://en.wikipedia.org/wiki/Bonaventure_des_P%C3%A9riers
Boniface Alexandre	http://en.wikipedia.org/wiki/Boniface_Alexandre
Bonnie Bedelia	http://en.wikipedia.org/wiki/Bonnie_Bedelia
Bonnie Blair	http://en.wikipedia.org/wiki/Bonnie_Blair
Bonnie Erbe	http://en.wikipedia.org/wiki/Bonnie_Erbe
Bonnie Franklin	http://en.wikipedia.org/wiki/Bonnie_Franklin
Bonnie Hunt	http://en.wikipedia.org/wiki/Bonnie_Hunt
Bonnie Parker	http://en.wikipedia.org/wiki/Bonnie_Parker
Bonnie Pointer	http://en.wikipedia.org/wiki/Bonnie_Pointer
Bonnie Raitt	http://en.wikipedia.org/wiki/Bonnie_Raitt
Bonnie Somerville	http://en.wikipedia.org/wiki/Bonnie_Somerville
Bonnie Tyler	http://en.wikipedia.org/wiki/Bonnie_Tyler
Bonny Lee Bakley	http://en.wikipedia.org/wiki/Bonny_Lee_Bakley
Boog Powell	http://en.wikipedia.org/wiki/Boog_Powell
Booker T	http://en.wikipedia.org/wiki/Booker_T._Jones
Booker T. Washington	http://en.wikipedia.org/wiki/Booker_T._Washington
Boomer Esiason	http://en.wikipedia.org/wiki/Boomer_Esiason
Booth Tarkington	http://en.wikipedia.org/wiki/Booth_Tarkington
Boots Randolph	http://en.wikipedia.org/wiki/Boots_Randolph
Bootsy Collins	http://en.wikipedia.org/wiki/Bootsy_Collins
Boris Altshuler	http://en.wikipedia.org/wiki/Boris_Altshuler
Boris Becker	http://en.wikipedia.org/wiki/Boris_Becker
Boris Blacher	http://en.wikipedia.org/wiki/Boris_Blacher
Boris Godunov	http://en.wikipedia.org/wiki/Boris_Godunov
Boris Karloff	http://en.wikipedia.org/wiki/Boris_Karloff
Boris Kodjoe	http://en.wikipedia.org/wiki/Boris_Kodjoe
Boris Pasternak	http://en.wikipedia.org/wiki/Boris_Pasternak
Boris Pickett	http://en.wikipedia.org/wiki/Boris_Pickett
Boris Spassky	http://en.wikipedia.org/wiki/Boris_Spassky
Boris Tadic	http://en.wikipedia.org/wiki/Boris_Tadi%C4%87
Boris Trajkovski	http://en.wikipedia.org/wiki/Boris_Trajkovski
Boris Vallejo	http://en.wikipedia.org/wiki/Boris_Vallejo
Boris Yeltsin	http://en.wikipedia.org/wiki/Boris_Yeltsin
Borislav Paravac	http://en.wikipedia.org/wiki/Borislav_Paravac
Borut Pahor	http://en.wikipedia.org/wiki/Borut_Pahor
Boss Tweed	http://en.wikipedia.org/wiki/Boss_Tweed
Bouasone Bouphavanh	http://en.wikipedia.org/wiki/Bouasone_Bouphavanh
Boungnang Vorachith	http://en.wikipedia.org/wiki/Boungnang_Vorachith
Bounty Killer	http://en.wikipedia.org/wiki/Bounty_Killer
Boutros Boutros-Ghali	http://en.wikipedia.org/wiki/Boutros_Boutros-Ghali
Bow Wow	http://en.wikipedia.org/wiki/Bow_Wow
Boxcar Willie	http://en.wikipedia.org/wiki/Boxcar_Willie
Boy George	http://en.wikipedia.org/wiki/Boy_George
Boyd Rice	http://en.wikipedia.org/wiki/Boyd_Rice
Boyko Borisov	http://en.wikipedia.org/wiki/Boyko_Borisov
Boz Burrell	http://en.wikipedia.org/wiki/Boz_Burrell
Boz Scaggs	http://en.wikipedia.org/wiki/Boz_Scaggs
Brad Bird	http://en.wikipedia.org/wiki/Brad_Bird
Brad Carson	http://en.wikipedia.org/wiki/Brad_Carson
Brad Davis	http://en.wikipedia.org/wiki/Brad_Davis_(actor)
Brad Delp	http://en.wikipedia.org/wiki/Brad_Delp
Brad Delson	http://en.wikipedia.org/wiki/Brad_Delson
Brad Dourif	http://en.wikipedia.org/wiki/Brad_Dourif
Brad Garrett	http://en.wikipedia.org/wiki/Brad_Garrett
Brad Henry	http://en.wikipedia.org/wiki/Brad_Henry
Brad Johnson	http://en.wikipedia.org/wiki/Brad_Johnson_%28American_football%29
Brad Miller	http://en.wikipedia.org/wiki/Brad_Miller_(congressman)
Brad Nowell	http://en.wikipedia.org/wiki/Brad_Nowell
Brad Paisley	http://en.wikipedia.org/wiki/Brad_Paisley
Brad Pitt	http://en.wikipedia.org/wiki/Brad_Pitt
Brad Renfro	http://en.wikipedia.org/wiki/Brad_Renfro
Brad Sherman	http://en.wikipedia.org/wiki/Brad_Sherman
Bradley Cooper	http://en.wikipedia.org/wiki/Bradley_Cooper
Bradley Whitford	http://en.wikipedia.org/wiki/Bradley_Whitford
Brady Anderson	http://en.wikipedia.org/wiki/Brady_Anderson
Bram Cohen	http://en.wikipedia.org/wiki/Bram_Cohen
Bram Stoker	http://en.wikipedia.org/wiki/Bram_Stoker
Brander Matthews	http://en.wikipedia.org/wiki/Brander_Matthews
Brandi Chastain	http://en.wikipedia.org/wiki/Brandi_Chastain
Brandon Albert	http://en.wikipedia.org/wiki/Brandon_Albert
Brandon Allen	http://en.wikipedia.org/wiki/Brandon_Allen
Brandon Boyd	http://en.wikipedia.org/wiki/Brandon_Boyd
Brandon Brooks	http://en.wikipedia.org/wiki/Brandon_Brooks_(actor)
Brandon Call	http://en.wikipedia.org/wiki/Brandon_Call
Brandon Cruz	http://en.wikipedia.org/wiki/Brandon_Cruz
Brandon De Wilde	http://en.wikipedia.org/wiki/Brandon_De_Wilde
Brandon DiCamillo	http://en.wikipedia.org/wiki/Brandon_DiCamillo
Brandon Flowers	http://en.wikipedia.org/wiki/Brandon_Flowers
Brandon Lee	http://en.wikipedia.org/wiki/Brandon_Lee
Brandon Lewis	http://en.wikipedia.org/wiki/Brandon_Lewis
Brandon Routh	http://en.wikipedia.org/wiki/Brandon_Routh
Brandy	http://en.wikipedia.org/wiki/Brandy_%28singer%29
Branford Marsalis	http://en.wikipedia.org/wiki/Branford_Marsalis
Brant Bjork	http://en.wikipedia.org/wiki/Brant_Bjork
Braxton Bragg	http://en.wikipedia.org/wiki/Braxton_Bragg
Breckin Meyer	http://en.wikipedia.org/wiki/Breckin_Meyer
Bree Sharp	http://en.wikipedia.org/wiki/Bree_Sharp
Brenda Bakke	http://en.wikipedia.org/wiki/Brenda_Bakke
Brenda Blethyn	http://en.wikipedia.org/wiki/Brenda_Blethyn
Brenda Fassie	http://en.wikipedia.org/wiki/Brenda_Fassie
Brenda Fricker	http://en.wikipedia.org/wiki/Brenda_Fricker
Brenda Holloway	http://en.wikipedia.org/wiki/Brenda_Holloway
Brenda K. Starr	http://en.wikipedia.org/wiki/Brenda_K._Starr
Brenda Lee	http://en.wikipedia.org/wiki/Brenda_Lee
Brenda Marshall	http://en.wikipedia.org/wiki/Brenda_Marshall
Brenda Song	http://en.wikipedia.org/wiki/Brenda_Song
Brenda Vaccaro	http://en.wikipedia.org/wiki/Brenda_Vaccaro
Brendan Behan	http://en.wikipedia.org/wiki/Brendan_Behan
Brendan Brazier	http://en.wikipedia.org/wiki/Brendan_Brazier
Brendan Eich	http://en.wikipedia.org/wiki/Brendan_Eich
Brendan Fehr	http://en.wikipedia.org/wiki/Brendan_Fehr
Brendan Fraser	http://en.wikipedia.org/wiki/Brendan_Fraser
Brendan T. Byrne	http://en.wikipedia.org/wiki/Brendan_T._Byrne
Brent Bozell	http://en.wikipedia.org/wiki/L._Brent_Bozell_III
Brent Briscoe	http://en.wikipedia.org/wiki/Brent_Briscoe
Brent Musburger	http://en.wikipedia.org/wiki/Brent_Musburger
Brent Scowcroft	http://en.wikipedia.org/wiki/Brent_Scowcroft
Brent Spiner	http://en.wikipedia.org/wiki/Brent_Spiner
Brent Wilkes	http://en.wikipedia.org/wiki/Brent_R._Wilkes
Bret Easton Ellis	http://en.wikipedia.org/wiki/Bret_Easton_Ellis
Bret Hart	http://en.wikipedia.org/wiki/Bret_Hart
Bret Harte	http://en.wikipedia.org/wiki/Bret_Harte
Bret Michaels	http://en.wikipedia.org/wiki/Bret_Michaels
Brett Anderson	http://en.wikipedia.org/wiki/Brett_Anderson
Brett Butler	http://en.wikipedia.org/wiki/Brett_Butler_(comedian)
Brett Favre	http://en.wikipedia.org/wiki/Brett_Favre
Brett Gurewitz	http://en.wikipedia.org/wiki/Brett_Gurewitz
Brett Guthrie	http://en.wikipedia.org/wiki/Brett_Guthrie
Brett Lee	http://en.wikipedia.org/wiki/Brett_Lee
Brett Ratner	http://en.wikipedia.org/wiki/Brett_Ratner
Brett Somers	http://en.wikipedia.org/wiki/Brett_Somers
Brian "Head" Welch	http://en.wikipedia.org/wiki/Brian_%22Head%22_Welch
Brian Aldiss	http://en.wikipedia.org/wiki/Brian_Aldiss
Brian Alford	http://en.wikipedia.org/wiki/Brian_Alford
Brian Allen	http://en.wikipedia.org/wiki/Brian_Allen_%28linebacker%29
Brian Anderson	http://en.wikipedia.org/wiki/Brian_Anderson_(skateboarder)
Brian Austin Green	http://en.wikipedia.org/wiki/Brian_Austin_Green
Brian Baird	http://en.wikipedia.org/wiki/Brian_Baird
Brian Bedford	http://en.wikipedia.org/wiki/Brian_Bedford
Brian Benben	http://en.wikipedia.org/wiki/Brian_Benben
Brian Bilbray	http://en.wikipedia.org/wiki/Brian_Bilbray
Brian Binley	http://en.wikipedia.org/wiki/Brian_Binley
Brian Blessed	http://en.wikipedia.org/wiki/Brian_Blessed
Brian Bloom	http://en.wikipedia.org/wiki/Brian_Bloom
Brian Boitano	http://en.wikipedia.org/wiki/Brian_Boitano
Brian Boru	http://en.wikipedia.org/wiki/Brian_Boru
Brian Bosworth	http://en.wikipedia.org/wiki/Brian_Bosworth
Brian Clough	http://en.wikipedia.org/wiki/Brian_Clough
Brian Cowen	http://en.wikipedia.org/wiki/Brian_Cowen
Brian Cox	http://en.wikipedia.org/wiki/Brian_Cox_(actor)
Brian D. Josephson	http://en.wikipedia.org/wiki/Brian_D._Josephson
Brian De Palma	http://en.wikipedia.org/wiki/Brian_De_Palma
Brian Dennehy	http://en.wikipedia.org/wiki/Brian_Dennehy
Brian Donlevy	http://en.wikipedia.org/wiki/Brian_Donlevy
Brian Donnelly	http://en.wikipedia.org/wiki/Brian_J._Donnelly
Brian Dougans	http://en.wikipedia.org/wiki/Brian_Dougans
Brian Doyle-Murray	http://en.wikipedia.org/wiki/Brian_Doyle-Murray
Brian Eno	http://en.wikipedia.org/wiki/Brian_Eno
Brian Epstein	http://en.wikipedia.org/wiki/Brian_Epstein
Brian France	http://en.wikipedia.org/wiki/Brian_France
Brian Friel	http://en.wikipedia.org/wiki/Brian_Friel
Brian Grazer	http://en.wikipedia.org/wiki/Brian_Grazer
Brian Greene	http://en.wikipedia.org/wiki/Brian_Greene
Brian Griese	http://en.wikipedia.org/wiki/Brian_Griese
Brian Helgeland	http://en.wikipedia.org/wiki/Brian_Helgeland
Brian Higgins	http://en.wikipedia.org/wiki/Brian_Higgins
Brian Hughes	http://en.wikipedia.org/wiki/Brian_Hughes_%28musician%29
Brian Johnson	http://en.wikipedia.org/wiki/Brian_Johnson
Brian Jones	http://en.wikipedia.org/wiki/Brian_Jones
Brian Keith	http://en.wikipedia.org/wiki/Brian_Keith
Brian Kernighan	http://en.wikipedia.org/wiki/Brian_Kernighan
Brian Kilmeade	http://en.wikipedia.org/wiki/Brian_Kilmeade
Brian Krause	http://en.wikipedia.org/wiki/Brian_Krause
Brian L. Roberts	http://en.wikipedia.org/wiki/Brian_L._Roberts
Brian Lamb	http://en.wikipedia.org/wiki/Brian_Lamb
Brian Lara	http://en.wikipedia.org/wiki/Brian_Lara
Brian Littrell	http://en.wikipedia.org/wiki/Brian_Littrell
Brian Maxwell	http://en.wikipedia.org/wiki/Brian_Maxwell
Brian May	http://en.wikipedia.org/wiki/Brian_May
Brian McKnight	http://en.wikipedia.org/wiki/Brian_McKnight
Brian Michael Bendis	http://en.wikipedia.org/wiki/Brian_Michael_Bendis
Brian Molko	http://en.wikipedia.org/wiki/Brian_Molko
Brian Moore	http://en.wikipedia.org/wiki/Brian_Moore_%28politician%29
Brian Mulroney	http://en.wikipedia.org/wiki/Brian_Mulroney
Brian Nichols	http://en.wikipedia.org/wiki/Brian_Nichols
Brian Posehn	http://en.wikipedia.org/wiki/Brian_Posehn
Brian Roberts	http://en.wikipedia.org/wiki/Brian_Roberts
Brian Ross	http://en.wikipedia.org/wiki/Brian_Ross_(journalist)
Brian Schweitzer	http://en.wikipedia.org/wiki/Brian_Schweitzer
Brian Setzer	http://en.wikipedia.org/wiki/Brian_Setzer
Brian Sibley	http://en.wikipedia.org/wiki/Brian_Sibley
Brian Sumner	http://en.wikipedia.org/wiki/Brian_Sumner
Brian Van Holt	http://en.wikipedia.org/wiki/Brian_Van_Holt
Brian Williams	http://en.wikipedia.org/wiki/Brian_Williams
Brian Wilson	http://en.wikipedia.org/wiki/Brian_Wilson
Bridget Fonda	http://en.wikipedia.org/wiki/Bridget_Fonda
Bridget Hall	http://en.wikipedia.org/wiki/Bridget_Hall
Bridget Moynahan	http://en.wikipedia.org/wiki/Bridget_Moynahan
Bridget Phillipson	http://en.wikipedia.org/wiki/Bridget_Phillipson
Bridgette Bardott	http://en.wikipedia.org/wiki/Brigit_Bardot
Bridgette Wilson	http://en.wikipedia.org/wiki/Bridgette_Wilson
Brigham Young	http://en.wikipedia.org/wiki/Brigham_Young
Brigid Brophy	http://en.wikipedia.org/wiki/Brigid_Brophy
Brigitte Bardot	http://en.wikipedia.org/wiki/Brigitte_Bardot
Brigitte Fontaine	http://en.wikipedia.org/wiki/Brigitte_Fontaine
Brigitte Mira	http://en.wikipedia.org/wiki/Brigitte_Mira
Brigitte Nielsen	http://en.wikipedia.org/wiki/Brigitte_Nielsen
Brini Maxwell	http://en.wikipedia.org/wiki/Brini_Maxwell
Brion Gysin	http://en.wikipedia.org/wiki/Brion_Gysin
Brion James	http://en.wikipedia.org/wiki/Brion_James
Brit Hume	http://en.wikipedia.org/wiki/Brit_Hume
Britney Spears	http://en.wikipedia.org/wiki/Britney_Spears
Britt Ekland	http://en.wikipedia.org/wiki/Britt_Ekland
Brittany Allen	http://en.wikipedia.org/wiki/Brittany_Allen
Brittany Daniel	http://en.wikipedia.org/wiki/Brittany_Daniel
Brittany Murphy	http://en.wikipedia.org/wiki/Brittany_Murphy
Brittany Snow	http://en.wikipedia.org/wiki/Brittany_Snow
Brock Adams	http://en.wikipedia.org/wiki/Brock_Adams
Brock Lesnar	http://en.wikipedia.org/wiki/Brock_Lesnar
Brock Peters	http://en.wikipedia.org/wiki/Brock_Peters
Brock Yates	http://en.wikipedia.org/wiki/Brock_Yates
Broderick Crawford	http://en.wikipedia.org/wiki/Broderick_Crawford
Brody Dalle	http://en.wikipedia.org/wiki/Brody_Dalle
Bronislaw Komorowski	http://en.wikipedia.org/wiki/Bronis%C5%82aw_Komorowski
Bronislaw Malinowski	http://en.wikipedia.org/wiki/Bronislaw_Malinowski
Bronson Alcott	http://en.wikipedia.org/wiki/Bronson_Alcott
Bronson Pinchot	http://en.wikipedia.org/wiki/Bronson_Pinchot
Brook Taylor	http://en.wikipedia.org/wiki/Brook_Taylor
Brooke Adams	http://en.wikipedia.org/wiki/Brooke_Adams_(actress)
Brooke Astor	http://en.wikipedia.org/wiki/Brooke_Astor
Brooke Burke	http://en.wikipedia.org/wiki/Brooke_Burke
Brooke Burns	http://en.wikipedia.org/wiki/Brooke_Burns
Brooke Langton	http://en.wikipedia.org/wiki/Brooke_Langton
Brooke Shields	http://en.wikipedia.org/wiki/Brooke_Shields
Brooke Valentine	http://en.wikipedia.org/wiki/Brooke_Shields
Brooks Adams	http://en.wikipedia.org/wiki/Brooks_Adams
Brooks Atkinson	http://en.wikipedia.org/wiki/Brooks_Atkinson
Brooks Newmark	http://en.wikipedia.org/wiki/Brooks_Newmark
Brooks Robinson	http://en.wikipedia.org/wiki/Brooks_Robinson
Bruce A. Morrison	http://en.wikipedia.org/wiki/Bruce_A._Morrison
Bruce Ackerman	http://en.wikipedia.org/wiki/Bruce_Ackerman
Bruce Allen	http://en.wikipedia.org/wiki/Bruce_Allen_%28American_football%29
Bruce Altman	http://en.wikipedia.org/wiki/Bruce_Altman
Bruce Babbitt	http://en.wikipedia.org/wiki/Bruce_Babbitt
Bruce Bagemihl	http://en.wikipedia.org/wiki/Bruce_Bagemihl
Bruce Bartlett	http://en.wikipedia.org/wiki/Bruce_Bartlett
Bruce Bennett	http://en.wikipedia.org/wiki/Bruce_Bennett
Bruce Beresford	http://en.wikipedia.org/wiki/Bruce_Beresford
Bruce Boxleitner	http://en.wikipedia.org/wiki/Bruce_Boxleitner
Bruce Braley	http://en.wikipedia.org/wiki/Bruce_Braley
Bruce Cabot	http://en.wikipedia.org/wiki/Bruce_Cabot
Bruce Campbell	http://en.wikipedia.org/wiki/Bruce_Campbell
Bruce Chatwin	http://en.wikipedia.org/wiki/Bruce_Chatwin
Bruce Cockburn	http://en.wikipedia.org/wiki/Bruce_Cockburn
Bruce Davidson	http://en.wikipedia.org/wiki/Bruce_Davidson_(photographer)
Bruce Davison	http://en.wikipedia.org/wiki/Bruce_Davison
Bruce Dern	http://en.wikipedia.org/wiki/Bruce_Dern
Bruce Dickinson	http://en.wikipedia.org/wiki/Bruce_Dickinson
Bruce E. Karatz	http://en.wikipedia.org/wiki/Bruce_Karatz
Bruce F. Vento	http://en.wikipedia.org/wiki/Bruce_F._Vento
Bruce Fein	http://en.wikipedia.org/wiki/Bruce_Fein
Bruce Golding	http://en.wikipedia.org/wiki/Bruce_Golding
Bruce Greenwood	http://en.wikipedia.org/wiki/Bruce_Greenwood
Bruce Haack	http://en.wikipedia.org/wiki/Bruce_Haack
Bruce Herschensohn	http://en.wikipedia.org/wiki/Bruce_Herschensohn
Bruce Hornsby	http://en.wikipedia.org/wiki/Bruce_Hornsby
Bruce Jenner	http://en.wikipedia.org/wiki/Bruce_Jenner
Bruce Lee	http://en.wikipedia.org/wiki/Bruce_Lee
Bruce Mahler	http://en.wikipedia.org/wiki/Bruce_Mahler
Bruce Marshall	http://en.wikipedia.org/wiki/Bruce_Marshall
Bruce McCulloch	http://en.wikipedia.org/wiki/Bruce_McCulloch
Bruce Merrifield	http://en.wikipedia.org/wiki/Bruce_Merrifield
Bruce Palmer	http://en.wikipedia.org/wiki/Bruce_Palmer
Bruce Ratner	http://en.wikipedia.org/wiki/Bruce_Ratner
Bruce Ritter	http://en.wikipedia.org/wiki/Bruce_Ritter
Bruce S. Gordon	http://en.wikipedia.org/wiki/Bruce_S._Gordon
Bruce Schneier	http://en.wikipedia.org/wiki/Bruce_Schneier
Bruce Shelley	http://en.wikipedia.org/wiki/Bruce_Shelley
Bruce Springsteen	http://en.wikipedia.org/wiki/Bruce_Springsteen
Bruce Sterling	http://en.wikipedia.org/wiki/Bruce_Sterling
Bruce Vento	http://en.wikipedia.org/wiki/Bruce_Vento
Bruce Vilanch	http://en.wikipedia.org/wiki/Bruce_Vilanch
Bruce Wasserstein	http://en.wikipedia.org/wiki/Bruce_Wasserstein
Bruce Willis	http://en.wikipedia.org/wiki/Bruce_Willis
Bruno Bettelheim	http://en.wikipedia.org/wiki/Bruno_Bettelheim
Bruno Frank	http://en.wikipedia.org/wiki/Bruno_Frank
Bruno Hauptmann	http://en.wikipedia.org/wiki/Bruno_Hauptmann
Bruno Kirby	http://en.wikipedia.org/wiki/Bruno_Kirby
Bruno Maderna	http://en.wikipedia.org/wiki/Bruno_Maderna
Bruno Nuytten	http://en.wikipedia.org/wiki/Bruno_Nuytten
Bryan Adams	http://en.wikipedia.org/wiki/Bryan_Adams
Bryan Brown	http://en.wikipedia.org/wiki/Bryan_Brown
Bryan Ferry	http://en.wikipedia.org/wiki/Bryan_Ferry
Bryan Forbes	http://en.wikipedia.org/wiki/Bryan_Forbes
Bryan Singer	http://en.wikipedia.org/wiki/Bryan_Singer
Bryant Gumbel	http://en.wikipedia.org/wiki/Bryant_Gumbel
Bryce Dallas Howard	http://en.wikipedia.org/wiki/Bryce_Dallas_Howard
Bryn Jones	http://en.wikipedia.org/wiki/Muslimgauze
Brynjar Aa	http://en.wikipedia.org/wiki/Brynjar_Aa
Bubba Baker	http://en.wikipedia.org/wiki/Bubba_Baker
Bubba Smith	http://en.wikipedia.org/wiki/Bubba_Smith
Buck 65	http://en.wikipedia.org/wiki/Buck_65
Buck Henry	http://en.wikipedia.org/wiki/Buck_Henry
Buck Jones	http://en.wikipedia.org/wiki/Buck_Jones
Buck McKeon	http://en.wikipedia.org/wiki/Buck_McKeon
Buck Owens	http://en.wikipedia.org/wiki/Buck_Owens
Bud Abbott	http://en.wikipedia.org/wiki/Bud_Abbott
Bud Cort	http://en.wikipedia.org/wiki/Bud_Cort
Bud Cramer	http://en.wikipedia.org/wiki/Bud_Cramer
Bud Lee	http://en.wikipedia.org/wiki/Bud_Lee
Bud McFarlane	http://en.wikipedia.org/wiki/Bud_McFarlane
Bud Powell	http://en.wikipedia.org/wiki/Bud_Powell
Bud Selig	http://en.wikipedia.org/wiki/Bud_Selig
Bud Shuster	http://en.wikipedia.org/wiki/Bud_Shuster
Bud Spencer	http://en.wikipedia.org/wiki/Bud_Spencer
Budd Boetticher	http://en.wikipedia.org/wiki/Budd_Boetticher
Budd Schulberg	http://en.wikipedia.org/wiki/Budd_Schulberg
Buddy Ebsen	http://en.wikipedia.org/wiki/Buddy_Ebsen
Buddy Guy	http://en.wikipedia.org/wiki/Buddy_Guy
Buddy Hackett	http://en.wikipedia.org/wiki/Buddy_Hackett
Buddy Holly	http://en.wikipedia.org/wiki/Buddy_Holly
Buddy MacKay	http://en.wikipedia.org/wiki/Buddy_MacKay
Buddy Rice	http://en.wikipedia.org/wiki/Buddy_Rice
Buddy Rich	http://en.wikipedia.org/wiki/Buddy_Rich
Buddy Rogers	http://en.wikipedia.org/wiki/Buddy_Rogers_%28wrestler%29
Buffalo Bill	http://en.wikipedia.org/wiki/Buffalo_Bill
Bug Hall	http://en.wikipedia.org/wiki/Bug_Hall
Bugsy Siegel	http://en.wikipedia.org/wiki/Bugsy_Siegel
Bulent Ecevit	http://en.wikipedia.org/wiki/Bulent_Ecevit
Bunny Berigan	http://en.wikipedia.org/wiki/Bunny_Berigan
Bunny DeBarge	http://en.wikipedia.org/wiki/Bunny_DeBarge
Bunny Lee	http://en.wikipedia.org/wiki/Bunny_Lee
Burgess Meredith	http://en.wikipedia.org/wiki/Burgess_Meredith
Burl Ives	http://en.wikipedia.org/wiki/Burl_Ives
Burt Bacharach	http://en.wikipedia.org/wiki/Burt_Bacharach
Burt Lancaster	http://en.wikipedia.org/wiki/Burt_Lancaster
Burt Reynolds	http://en.wikipedia.org/wiki/Burt_Reynolds
Burt Rutan	http://en.wikipedia.org/wiki/Burt_Rutan
Burt Ward	http://en.wikipedia.org/wiki/Burt_Ward
Burt Young	http://en.wikipedia.org/wiki/Burt_Young
Burton Richardson	http://en.wikipedia.org/wiki/Burton_Richardson
Burton Richter	http://en.wikipedia.org/wiki/Burton_Richter
Busby Berkeley	http://en.wikipedia.org/wiki/Busby_Berkeley
Busta Rhymes	http://en.wikipedia.org/wiki/Busta_Rhymes
Buster Crabbe	http://en.wikipedia.org/wiki/Buster_Crabbe
Buster Keaton	http://en.wikipedia.org/wiki/Buster_Keaton
Butch Otter	http://en.wikipedia.org/wiki/Butch_Otter
Butch Patrick	http://en.wikipedia.org/wiki/Butch_Patrick
Butch Vig	http://en.wikipedia.org/wiki/Butch_Vig
Butler Derrick	http://en.wikipedia.org/wiki/Butler_Derrick
Butterfly McQueen	http://en.wikipedia.org/wiki/Butterfly_McQueen
Button Gwinnett	http://en.wikipedia.org/wiki/Button_Gwinnett
Buzz Aldrin	http://en.wikipedia.org/wiki/Buzz_Aldrin
Buzz Osborne	http://en.wikipedia.org/wiki/Buzz_Osborne
Byron Allen	http://en.wikipedia.org/wiki/Byron_Allen
Byron Dorgan	http://en.wikipedia.org/wiki/Byron_Dorgan
Byron Grote	http://en.wikipedia.org/wiki/Byron_Grote
Byron L. Dorgan	http://en.wikipedia.org/wiki/Byron_L._Dorgan
Byron Nelson	http://en.wikipedia.org/wiki/Byron_Nelson
Byron White	http://en.wikipedia.org/wiki/Byron_White
Byron York	http://en.wikipedia.org/wiki/Byron_York
C. Aubrey Smith	http://en.wikipedia.org/wiki/C._Aubrey_Smith
C. Boyden Gray	http://en.wikipedia.org/wiki/C._Boyden_Gray
C. Delores Tucker	http://en.wikipedia.org/wiki/C._Delores_Tucker
C. Douglas Dillon	http://en.wikipedia.org/wiki/C._Douglas_Dillon
C. Everett Koop	http://en.wikipedia.org/wiki/C._Everett_Koop
C. Hartley Grattan	http://en.wikipedia.org/wiki/C._Hartley_Grattan
C. J. Cherryh	http://en.wikipedia.org/wiki/C._J._Cherryh
C. K. Williams	http://en.wikipedia.org/wiki/C._K._Williams
C. M. Kornbluth	http://en.wikipedia.org/wiki/C._M._Kornbluth
C. Martin Croker	http://en.wikipedia.org/wiki/C._Martin_Croker
C. Michael Armstrong	http://en.wikipedia.org/wiki/C._Michael_Armstrong
C. P. Snow	http://en.wikipedia.org/wiki/C._P._Snow
C. S. Forester	http://en.wikipedia.org/wiki/C._S._Forester
C. S. Lewis	http://en.wikipedia.org/wiki/C._S._Lewis
C. T. R. Wilson	http://en.wikipedia.org/wiki/C._T._R._Wilson
C. Thomas Howell	http://en.wikipedia.org/wiki/C._Thomas_Howell
C. Vann Woodward	http://en.wikipedia.org/wiki/C._Vann_Woodward
C. William Verity	http://en.wikipedia.org/wiki/C._William_Verity
C. Wright Mills	http://en.wikipedia.org/wiki/C._Wright_Mills
C.C. DeVille	http://en.wikipedia.org/wiki/C.C._DeVille
C.W. Bill Young	http://en.wikipedia.org/wiki/C.W._Bill_Young
Cab Calloway	http://en.wikipedia.org/wiki/Cab_Calloway
Cadwallader Colden Washburn	http://en.wikipedia.org/wiki/Cadwallader_Colden_Washburn
Caesar Augustus	http://en.wikipedia.org/wiki/Caesar_Augustus
Caetano Veloso	http://en.wikipedia.org/wiki/Caetano_Veloso
Caitlin Flanagan	http://en.wikipedia.org/wiki/Caitlin_Flanagan
Cal Dooley	http://en.wikipedia.org/wiki/Cal_Dooley
Cal Ripken	http://en.wikipedia.org/wiki/Cal_Ripken
Cal Thomas	http://en.wikipedia.org/wiki/Cal_Thomas
Cal Tjader	http://en.wikipedia.org/wiki/Cal_Tjader
Cal Worthington	http://en.wikipedia.org/wiki/Cal_Worthington
Calamity Jane	http://en.wikipedia.org/wiki/Calamity_Jane
Cale Yarborough	http://en.wikipedia.org/wiki/Cale_Yarborough
Caleb Cushing	http://en.wikipedia.org/wiki/Caleb_Cushing
Calin Popescu-Tariceanu	http://en.wikipedia.org/wiki/Calin_Popescu-Tariceanu
Calista Flockhart	http://en.wikipedia.org/wiki/Calista_Flockhart
Calisto Tanzi	http://en.wikipedia.org/wiki/Calisto_Tanzi
Calvert DeForest	http://en.wikipedia.org/wiki/Calvert_DeForest
Calvin Coolidge	http://en.wikipedia.org/wiki/Calvin_Coolidge
Calvin Klein	http://en.wikipedia.org/wiki/Calvin_Klein_(fashion_designer)
Calvin Murphy	http://en.wikipedia.org/wiki/Calvin_Murphy
Calvin Trillin	http://en.wikipedia.org/wiki/Calvin_Trillin
Cameron Crowe	http://en.wikipedia.org/wiki/Cameron_Crowe
Cameron Diaz	http://en.wikipedia.org/wiki/Cameron_Diaz
Cameron Dye	http://en.wikipedia.org/wiki/Cameron_Dye
Cameron Kerry	http://en.wikipedia.org/wiki/Cameron_Kerry
Cameron Mitchell	http://en.wikipedia.org/wiki/Cameron_Mitchell_(actor)
Camilla Parker Bowles	http://en.wikipedia.org/wiki/Camilla_Parker_Bowles
Camille Claudel	http://en.wikipedia.org/wiki/Camille_Claudel
Camille Corot	http://en.wikipedia.org/wiki/Camille_Corot
Camille Desmoulins	http://en.wikipedia.org/wiki/Camille_Desmoulins
Camille Paglia	http://en.wikipedia.org/wiki/Camille_Paglia
Camille Pissarro	http://en.wikipedia.org/wiki/Camille_Pissarro
Camille Saint-Sa�ns	http://en.wikipedia.org/wiki/Camille_Saint-Sa%C3%Abns
Camillo Benso di Cavour	http://en.wikipedia.org/wiki/Camillo_Benso_di_Cavour
Camilo Jos� Cela	http://en.wikipedia.org/wiki/Camilo_Jos%C3%A9_Cela
Campbell Brown	http://en.wikipedia.org/wiki/Campbell_Brown
Campbell Scott	http://en.wikipedia.org/wiki/Campbell_Scott
Camryn Manheim	http://en.wikipedia.org/wiki/Camryn_Manheim
Candace Allen	http://en.wikipedia.org/wiki/Candace_Allen
Candace Bergan	http://en.wikipedia.org/wiki/Candice_Bergen
Candace Bushnell	http://en.wikipedia.org/wiki/Candace_Bushnell
Candace Cameron	http://en.wikipedia.org/wiki/Candace_Cameron
Candice Bergen	http://en.wikipedia.org/wiki/Candice_Bergen
Candice Miller	http://en.wikipedia.org/wiki/Candice_Miller
Candy Barr	http://en.wikipedia.org/wiki/Candy_Barr
Candy Crowley	http://en.wikipedia.org/wiki/Candy_Crowley
Cannonball Adderley	http://en.wikipedia.org/wiki/Cannonball_Adderley
Caprice Bourret	http://en.wikipedia.org/wiki/Caprice_Bourret
Captain Beefheart	http://en.wikipedia.org/wiki/Captain_Beefheart
Captain Crunch	http://en.wikipedia.org/wiki/John_Draper
Captain Kangaroo	http://en.wikipedia.org/wiki/Captain_Kangaroo
Captain Lou Albano	http://en.wikipedia.org/wiki/Captain_Lou_Albano
Captain Sensible	http://en.wikipedia.org/wiki/Captain_Sensible
Cardinal Richelieu	http://en.wikipedia.org/wiki/Cardinal_Richelieu
Cardiss Collins	http://en.wikipedia.org/wiki/Cardiss_Collins
Carey Hart	http://en.wikipedia.org/wiki/Carey_Hart
Carey Lowell	http://en.wikipedia.org/wiki/Carey_Lowell
Carey McWilliams	http://en.wikipedia.org/wiki/Carey_McWilliams_(journalist)
Carey Means	http://en.wikipedia.org/wiki/Carey_Means
Carl Adams	http://en.wikipedia.org/wiki/Carl_Adams
Carl Akeley	http://en.wikipedia.org/wiki/Carl_Akeley
Carl Allen	http://en.wikipedia.org/wiki/Carl_Allen_%28American_football%29
Carl B. Albert	http://en.wikipedia.org/wiki/Carl_B._Albert
Carl Bar�t	http://en.wikipedia.org/wiki/Carl_Bar%C3%A2t
Carl Becker	http://en.wikipedia.org/wiki/Carl_Becker_%28general%29
Carl Bernstein	http://en.wikipedia.org/wiki/Carl_Bernstein
Carl Betz	http://en.wikipedia.org/wiki/Carl_Betz
Carl Bosch	http://en.wikipedia.org/wiki/Carl_Bosch
Carl C. Perkins	http://en.wikipedia.org/wiki/Carl_C._Perkins
Carl Cameron	http://en.wikipedia.org/wiki/Carl_Cameron
Carl Czerny	http://en.wikipedia.org/wiki/Carl_Czerny
Carl D. Pursell	http://en.wikipedia.org/wiki/Carl_D._Pursell
Carl David Anderson	http://en.wikipedia.org/wiki/Carl_David_Anderson
Carl E. Wieman	http://en.wikipedia.org/wiki/Carl_E._Wieman
Carl Friedrich Gauss	http://en.wikipedia.org/wiki/Carl_Friedrich_Gauss
Carl Goerdeler	http://en.wikipedia.org/wiki/Carl_Goerdeler
Carl Gustaf Emil Mannerheim	http://en.wikipedia.org/wiki/Carl_Gustaf_Emil_Mannerheim
Carl Gustaf, Count Tessin	http://en.wikipedia.org/wiki/Carl_Gustaf_Tessin
Carl Hiaasen	http://en.wikipedia.org/wiki/Carl_Hiaasen
Carl Hubbell	http://en.wikipedia.org/wiki/Carl_Hubbell
Carl Icahn	http://en.wikipedia.org/wiki/Carl_Icahn
Carl Jung	http://en.wikipedia.org/wiki/Carl_Jung
Carl Karcher	http://en.wikipedia.org/wiki/Carl_Karcher
Carl Kasell	http://en.wikipedia.org/wiki/Carl_Kasell
Carl Levin	http://en.wikipedia.org/wiki/Carl_Levin
Carl Lewis	http://en.wikipedia.org/wiki/Carl_Lewis
Carl Loewe	http://en.wikipedia.org/wiki/Carl_Loewe
Carl Malamud	http://en.wikipedia.org/wiki/Carl_Malamud
Carl Maria von Weber	http://en.wikipedia.org/wiki/Carl_Maria_von_Weber
Carl Nielsen	http://en.wikipedia.org/wiki/Carl_Nielsen
Carl Orff	http://en.wikipedia.org/wiki/Carl_Orff
Carl Palmer	http://en.wikipedia.org/wiki/Carl_Palmer
Carl Perkins	http://en.wikipedia.org/wiki/Carl_Perkins
Carl Pope	http://en.wikipedia.org/wiki/Carl_Pope
Carl Reiner	http://en.wikipedia.org/wiki/Carl_Reiner
Carl Remigius Fresenius	http://en.wikipedia.org/wiki/Carl_Remigius_Fresenius
Carl Rowan	http://en.wikipedia.org/wiki/Carl_Rowan
Carl Sagan	http://en.wikipedia.org/wiki/Carl_Sagan
Carl Sandburg	http://en.wikipedia.org/wiki/Carl_Sandburg
Carl Stalling	http://en.wikipedia.org/wiki/Carl_Stalling
Carl Switzer	http://en.wikipedia.org/wiki/Carl_Switzer
Carl Theodor Dreyer	http://en.wikipedia.org/wiki/Carl_Switzer
Carl Van Doren	http://en.wikipedia.org/wiki/Carl_Van_Doren
Carl Van Vechten	http://en.wikipedia.org/wiki/Carl_Van_Vechten
Carl von Clausewitz	http://en.wikipedia.org/wiki/Carl_von_Clausewitz
Carl von Cosel	http://en.wikipedia.org/wiki/Carl_von_Cosel
Carl von Ossietzky	http://en.wikipedia.orghttp://en.wikipedia.org/wiki/Carl_von_Ossietzky
Carl Weathers	http://en.wikipedia.org/wiki/Carl_Weathers
Carl Wilhelm Scheele	http://en.wikipedia.org/wiki/Carl_Wilhelm_Scheele
Carl Wilson	http://en.wikipedia.org/wiki/Carl_Wilson
Carl XVI Gustaf	http://en.wikipedia.org/wiki/Carl_XVI_Gustaf
Carl Yastrzemski	http://en.wikipedia.org/wiki/Carl_Yastrzemski
Carla Bley	http://en.wikipedia.org/wiki/Carla_Bley
Carla Gugino	http://en.wikipedia.org/wiki/Carla_Gugino
Carl-Henric Svanberg	http://en.wikipedia.org/wiki/Carl-Henric_Svanberg
Carlie Brucia	http://en.wikipedia.org/w/index.php?title=Carlie_Brucia
Carlo Allen	http://en.wikipedia.org/wiki/Carlos_Allen
Carlo Azeglio Ciampi	http://en.wikipedia.org/wiki/Carlo_Azeglio_Ciampi
Carlo Crivelli	http://en.wikipedia.org/wiki/Carlo_Crivelli
Carlo Denina	http://en.wikipedia.org/wiki/Carlo_Denina
Carlo Gambino	http://en.wikipedia.org/wiki/Carlo_Gambino
Carlo Goldoni	http://en.wikipedia.org/wiki/Carlo_Goldoni
Carlo Passaglia	http://en.wikipedia.org/wiki/Carlo_Passaglia
Carlo Perez Allen	http://en.wikipedia.org/wiki/Carlos_Allen
Carlo Ponti	http://en.wikipedia.org/wiki/Carlo_Ponti
Carlo Rubbia	http://en.wikipedia.org/wiki/Carlo_Rubbia
Carlos Alazraqui	http://en.wikipedia.org/wiki/Carlos_Alazraqui
Carlos Allen	http://en.wikipedia.org/wiki/Carlos_Allen
Carlos Alomar	http://en.wikipedia.org/wiki/Carlos_Alomar
Carlos Castaneda	http://en.wikipedia.org/wiki/Carlos_Castaneda
Carlos Ch�vez	http://en.wikipedia.org/wiki/Carlos_Ch%C3%A1vez
Carlos de Sig�enza y G�ngora	http://en.wikipedia.org/wiki/Carlos_de_Sig%C3%BCenza_y_G%C3%B3ngora
Carlos de Sig�enza y G�ngora	http://en.wikipedia.org/wiki/Carlos_de_Sig%C3%BCenza_y_G%C3%B3ngora
Carlos Filipe Ximenes Belo	http://en.wikipedia.org/wiki/Carlos_Filipe_Ximenes_Belo
Carlos Fuentes	http://en.wikipedia.org/wiki/Carlos_Fuentes
Carlos Gomes J�nior	http://en.wikipedia.org/wiki/Carlos_Gomes_J%C3%Banior
Carlos Gutierrez	http://en.wikipedia.org/wiki/Carlos_Gutierrez
Carlos J. Moorhead	http://en.wikipedia.org/wiki/Carlos_J._Moorhead
Carlos Mencia	http://en.wikipedia.org/wiki/Carlos_Mencia
Carlos Menem	http://en.wikipedia.org/wiki/Carlos_Menem
Carlos Mesa	http://en.wikipedia.org/wiki/Carlos_Mesa
Carlos P. Garcia	http://en.wikipedia.org/wiki/Carlos_P._Garcia
Carlos Ponce	http://en.wikipedia.org/wiki/Carlos_Ponce
Carlos Saavedra Lamas	http://en.wikipedia.org/wiki/Carlos_Saavedra_Lamas
Carlos Salinas	http://en.wikipedia.org/wiki/Carlos_Salinas
Carlos Santana	http://en.wikipedia.org/wiki/Carlos_Santana
Carlos Slim Helu	http://en.wikipedia.org/wiki/Carlos_Slim_Helu
Carlos T�vez	http://en.wikipedia.org/wiki/Carlos_T%C3%A9vez
Carlos the Jackal	http://en.wikipedia.org/wiki/Carlos_the_Jackal
Carlton Fisk	http://en.wikipedia.org/wiki/Carlton_Fisk
Carly Fiorina	http://en.wikipedia.org/wiki/Carly_Fiorina
Carly Pope	http://en.wikipedia.org/wiki/Carly_Pope
Carly Simon	http://en.wikipedia.org/wiki/Carly_Simon
Carmelo Anthony	http://en.wikipedia.org/wiki/Carmelo_Anthony
Carmen Alvarez	http://en.wikipedia.org/wiki/Carmen_Julia_%C3%81lvarez
Carmen Electra	http://en.wikipedia.org/wiki/Carmen_Electra
Carmen Kass	http://en.wikipedia.org/wiki/Carmen_Kass
Carmen Miranda	http://en.wikipedia.org/wiki/Carmen_Miranda
Carmine Appice	http://en.wikipedia.org/wiki/Carmine_Appice
Carmine De Sapio	http://en.wikipedia.org/wiki/Carmine_De_Sapio
Carnie Wilson	http://en.wikipedia.org/wiki/Carnie_Wilson
Carol Allen	http://en.wikipedia.org/wiki/Carol_Allen
Carol Alt	http://en.wikipedia.org/wiki/Carol_Alt
Carol Ann Duffy	http://en.wikipedia.org/wiki/Carol_Ann_Duffy
Carol Bruce	http://en.wikipedia.org/wiki/Carol_Bruce
Carol Burnett	http://en.wikipedia.org/wiki/Carol_Burnett
Carol Channing	http://en.wikipedia.org/wiki/Carol_Channing
Carol Doda	http://en.wikipedia.org/wiki/Carol_Doda
Carol Gilligan	http://en.wikipedia.org/wiki/Carol_Gilligan
Carol Kane	http://en.wikipedia.org/wiki/Carol_Kane
Carol Leifer	http://en.wikipedia.org/wiki/Carol_Leifer
Carol Lynley	http://en.wikipedia.org/wiki/Carol_Lynley
Carol M. Browner	http://en.wikipedia.org/wiki/Carol_M._Browner
Carol Moseley Braun	http://en.wikipedia.org/wiki/Carol_Moseley_Braun
Carol Reed	http://en.wikipedia.org/wiki/Carol_Reed
Carol Shea-Porter	http://en.wikipedia.org/wiki/Carol_Shea-Porter
Carol Shields	http://en.wikipedia.org/wiki/Carol_Shields
Carol Wayne	http://en.wikipedia.org/wiki/Carol_Wayne
Carole King	http://en.wikipedia.org/wiki/Carole_King
Carole Landis	http://en.wikipedia.org/wiki/Carole_Landis
Carole Lombard	http://en.wikipedia.org/wiki/Carole_Lombard
Caroline B. Cooney	http://en.wikipedia.org/wiki/Caroline_B._Cooney
Caroline Dinenage	http://en.wikipedia.org/wiki/Caroline_Dinenage
Caroline Flint	http://en.wikipedia.org/wiki/Caroline_Flint
Caroline Herschel	http://en.wikipedia.org/wiki/Caroline_Herschel
Caroline Kennedy	http://en.wikipedia.org/wiki/Caroline_Kennedy
Caroline Lucas	http://en.wikipedia.org/wiki/Caroline_Lucas
Caroline Nokes	http://en.wikipedia.org/wiki/Caroline_Nokes
Caroline Spelman	http://en.wikipedia.org/wiki/Caroline_Spelman
Caroll Spinney	http://en.wikipedia.org/wiki/Caroll_Spinney
Carolus Linnaeus	http://en.wikipedia.org/wiki/Carolus_Linnaeus
Carolyn Cassady	http://en.wikipedia.org/wiki/Carolyn_Cassady
Carolyn Forché	http://en.wikipedia.org/wiki/Carolyn_Forch%C3%A9
Carolyn Heilbrun	http://en.wikipedia.org/wiki/Carolyn_Heilbrun
Carolyn Jones	http://en.wikipedia.org/wiki/Carolyn_Jones
Carolyn Kilpatrick	http://en.wikipedia.org/wiki/Carolyn_Kilpatrick
Carolyn Kizer	http://en.wikipedia.org/wiki/Carolyn_Kizer
Carolyn Maloney	http://en.wikipedia.org/wiki/Carolyn_Maloney
Carolyn McCarthy	http://en.wikipedia.org/wiki/Carolyn_McCarthy
Carolyn Meinel	http://en.wikipedia.org/wiki/Carolyn_Meinel
Caron Keating	http://en.wikipedia.org/wiki/Caron_Keating
Carre Otis	http://en.wikipedia.org/wiki/Carre_Otis
Carr� Otis	http://en.wikipedia.org/wiki/Carr%C3%A9_Otis
Carrie Allen	http://en.wikipedia.org/wiki/Carrie_Allen#Carrie_Allen
Carrie Fisher	http://en.wikipedia.org/wiki/Carrie_Fisher
Carrie Henn	http://en.wikipedia.org/wiki/Carrie_Henn
Carrie Nation	http://en.wikipedia.org/wiki/Carrie_Nation
Carrie P. Meek	http://en.wikipedia.org/wiki/Carrie_P._Meek
Carrie Snodgress	http://en.wikipedia.org/wiki/Carrie_Snodgress
Carrie Underwood	http://en.wikipedia.org/wiki/Carrie_Underwood
Carrie-Anne Moss	http://en.wikipedia.org/wiki/Carrie-Anne_Moss
Carroll A. Campbell, Jr.	http://en.wikipedia.org/wiki/Carroll_A._Campbell%2C_Jr.
Carroll Baker	http://en.wikipedia.org/wiki/Carroll_Baker
Carroll Campbell	http://en.wikipedia.org/wiki/Carroll_Campbell
Carroll Hubbard, Jr.	http://en.wikipedia.org/wiki/Carroll_Hubbard%2C_Jr.
Carroll O'Connor	http://en.wikipedia.org/wiki/Carroll_O%27Connor
Carroll Shelby	http://en.wikipedia.org/wiki/Carroll_Shelby
Carrot Top	http://en.wikipedia.org/wiki/Carrot_Top
Carson Daly	http://en.wikipedia.org/wiki/Carson_Daly
Carson Kressley	http://en.wikipedia.org/wiki/Carson_Kressley
Carson McCullers	http://en.wikipedia.org/wiki/Carson_McCullers
Carsten Nicolai	http://en.wikipedia.org/wiki/Carsten_Nicolai
Carter Burwell	http://en.wikipedia.org/wiki/Carter_Burwell
Carter Oosterhouse	http://en.wikipedia.org/wiki/Carter_Oosterhouse
Carter T. Barron	http://en.wikipedia.org/w/index.php?title=Carter_T._Barron
Cary Elwes	http://en.wikipedia.org/wiki/Cary_Elwes
Cary Grant	http://en.wikipedia.org/wiki/Cary_Grant
Cary Stayner	http://en.wikipedia.org/wiki/Cary_Stayner
Caryl Churchill	http://en.wikipedia.org/wiki/Caryl_Churchill
Caryl Phillips	http://en.wikipedia.org/wiki/Caryl_Phillips
Casey Affleck	http://en.wikipedia.org/wiki/Casey_Affleck
Casey Kasem	http://en.wikipedia.org/wiki/Casey_Kasem
Casey Stengel	http://en.wikipedia.org/wiki/Casey_Stengel
Casimir Delavigne	http://en.wikipedia.org/wiki/Casimir_Delavigne
Casimir III	http://en.wikipedia.org/wiki/Casimir_III_of_Poland
Casimir IV	http://en.wikipedia.org/wiki/Casimir_IV_Jagiellon
Casimir Pulaski	http://en.wikipedia.org/wiki/Casimir_Pulaski
Caspar David Friedrich	http://en.wikipedia.org/wiki/Caspar_David_Friedrich
Caspar Weinberger	http://en.wikipedia.org/wiki/Caspar_Weinberger
Casper Van Dien	http://en.wikipedia.org/wiki/Casper_Van_Dien
Cass Ballenger	http://en.wikipedia.org/wiki/Cass_Ballenger
Cass Sunstein	http://en.wikipedia.org/wiki/Cass_Sunstein
Cassandra Wilson	http://en.wikipedia.org/wiki/Cassandra_Wilson
Cassius Marcellus Clay	http://en.wikipedia.org/wiki/Cassius_Marcellus_Clay_%281810%E2%80%931903%29
Cassius Marcellus Coolidge	http://en.wikipedia.org/wiki/Cassius_Marcellus_Coolidge
Cat Stevens	http://en.wikipedia.org/wiki/Cat_Stevens
Cate Blanchett	http://en.wikipedia.org/wiki/Cate_Blanchett
Catfish Hunter	http://en.wikipedia.org/wiki/Catfish_Hunter
Cath Carroll	http://en.wikipedia.org/wiki/Cath_Carroll
Catharine MacKinnon	http://en.wikipedia.org/wiki/Catharine_MacKinnon
Catherine Bach	http://en.wikipedia.org/wiki/Catherine_Bach
Catherine Bell	http://en.wikipedia.org/wiki/Catherine_Bell
Catherine Crier	http://en.wikipedia.org/wiki/Catherine_Crier
Catherine de Medici	http://en.wikipedia.org/wiki/Catherine_de_Medici
Catherine Deneuve	http://en.wikipedia.org/wiki/Catherine_Deneuve
Catherine Hicks	http://en.wikipedia.org/wiki/Catherine_Hicks
Catherine Howard	http://en.wikipedia.org/wiki/Catherine_Howard
Catherine I	http://en.wikipedia.org/wiki/Catherine_I
Catherine Keener	http://en.wikipedia.org/wiki/Catherine_Keener
Catherine McCormack	http://en.wikipedia.org/wiki/Catherine_McCormack
Catherine McKinnell	http://en.wikipedia.org/wiki/Catherine_McKinnell
Catherine of Aragon	http://en.wikipedia.org/wiki/Catherine_of_Aragon
Catherine of Braganza	http://en.wikipedia.org/wiki/Catherine_of_Braganza
Catherine of Valois	http://en.wikipedia.org/wiki/Catherine_of_Valois
Catherine O'Hara	http://en.wikipedia.org/wiki/Catherine_O%27Hara
Catherine Oxenberg	http://en.wikipedia.org/wiki/Catherine_Oxenberg
Catherine Parr	http://en.wikipedia.org/wiki/Catherine_Parr
Catherine S. Long	http://en.wikipedia.org/wiki/Catherine_S._Long
Catherine Swynford	http://en.wikipedia.org/wiki/Catherine_Swynford
Catherine the Great	http://en.wikipedia.org/wiki/Catherine_the_Great
Catherine Zeta-Jones	http://en.wikipedia.org/wiki/Catherine_Zeta-Jones
Cathy Dennis	http://en.wikipedia.org/wiki/Cathy_Dennis
Cathy Guisewite	http://en.wikipedia.org/wiki/Cathy_Guisewite
Cathy Jamieson	http://en.wikipedia.org/wiki/Cathy_Jamieson
Cathy Lee Crosby	http://en.wikipedia.org/wiki/Cathy_Lee_Crosby
Cathy McMorris	http://en.wikipedia.org/wiki/Cathy_McMorris
Cathy Moriarty	http://en.wikipedia.org/wiki/Cathy_Moriarty
Cathy Rigby	http://en.wikipedia.org/wiki/Cathy_Rigby
Cato the Elder	http://en.wikipedia.org/wiki/Cato_the_Elder
Cato the Younger	http://en.wikipedia.org/wiki/Cato_the_Younger
CCH Pounder	http://en.wikipedia.org/wiki/CCH_Pounder
Cecil Adams	http://en.wikipedia.org/wiki/Cecil_Adams
Cecil B. DeMille	http://en.wikipedia.org/wiki/Cecil_B._DeMille
Cecil D. Andrus	http://en.wikipedia.org/wiki/Cecil_D._Andrus
Cecil Day-Lewis	http://en.wikipedia.org/wiki/Cecil_Day-Lewis
Cecil Fielder	http://en.wikipedia.org/wiki/Cecil_Fielder
Cecil Heftel	http://en.wikipedia.org/wiki/Cecil_Heftel
Cecil Kellaway	http://en.wikipedia.org/wiki/Cecil_Kellaway
Cecil Powell	http://en.wikipedia.org/wiki/Cecil_Powell
Cecil Rhodes	http://en.wikipedia.org/wiki/Cecil_Rhodes
Cecil Taylor	http://en.wikipedia.org/wiki/Cecil_Taylor
Cecile Dionne	http://en.wikipedia.org/wiki/Cecile_Dionne
Cecilia Parker	http://en.wikipedia.org/wiki/Cecilia_Parker
Cedric Hardwicke	http://en.wikipedia.org/wiki/Cedric_Hardwicke
Cedric the Entertainer	http://en.wikipedia.org/wiki/Cedric_the_Entertainer
Cedric Yarbrough	http://en.wikipedia.org/wiki/Cedric_Yarbrough
Cele Abba	http://en.wikipedia.org/wiki/Cele_Abba
Celeste Holm	http://en.wikipedia.org/wiki/Celeste_Holm
Celia Cruz	http://en.wikipedia.org/wiki/Celia_Cruz
Celia Johnson	http://en.wikipedia.org/wiki/Celia_Johnson
Celine Dion	http://en.wikipedia.org/wiki/Celine_Dion
Cellou Dalein Diallo	http://en.wikipedia.org/wiki/Cellou_Dalein_Diallo
Cesar Amigo	http://en.wikipedia.org/wiki/Cesar_Amigo
Cesar Chavez	http://en.wikipedia.org/wiki/Cesar_Chavez
C�sar Franck	http://en.wikipedia.org/wiki/C%C3%A9sar_Franck
Cesar Romero	http://en.wikipedia.org/wiki/Cesar_Romero
Cesare Borgia	http://en.wikipedia.org/wiki/Cesare_Borgia
Cesare Pavese	http://en.wikipedia.org/wiki/Cesare_Pavese
cEvin Key	http://en.wikipedia.org/wiki/cEvin_Key
Chad Allen	http://en.wikipedia.org/wiki/Chad_Allen_(actor)
Chad Everett	http://en.wikipedia.org/wiki/Chad_Everett
Chad Hugo	http://en.wikipedia.org/wiki/Chad_Hugo
Chad Kroeger	http://en.wikipedia.org/wiki/Chad_Kroeger
Chad Lowe	http://en.wikipedia.org/wiki/Chad_Lowe
Chad Michael Murray	http://en.wikipedia.org/wiki/Chad_Michael_Murray
Chad Smith	http://en.wikipedia.org/wiki/Chad_Smith
Chae An	http://en.wikipedia.org/wiki/Chae_An
Chaim Herzog	http://en.wikipedia.org/wiki/Chaim_Herzog
Chaim Potok	http://en.wikipedia.org/wiki/Chaim_Potok
Chaim Soutine	http://en.wikipedia.org/wiki/Chaim_Soutine
Chaim Weizmann	http://en.wikipedia.org/wiki/Chaim_Weizmann
Chaka Fattah	http://en.wikipedia.org/wiki/Chaka_Fattah
Chaka Khan	http://en.wikipedia.org/wiki/Chaka_Khan
Chalino Sanchez	http://en.wikipedia.org/wiki/Chalino_Sanchez
Chalmers P. Wylie	http://en.wikipedia.org/wiki/Chalmers_P._Wylie
Chaminda Vaas	http://en.wikipedia.org/wiki/Chaminda_Vaas
Chan Marshall	http://en.wikipedia.org/wiki/Chan_Marshall
Chan Romero	http://en.wikipedia.org/wiki/Chan_Romero
Chandler Brossard	http://en.wikipedia.org/wiki/Chandler_Brossard
Chandra Levy	http://en.wikipedia.org/wiki/Chandra_Levy
Chandrasekhara Venkata Raman	http://en.wikipedia.org/wiki/Chandrasekhara_Venkata_Raman
Channing Tatum	http://en.wikipedia.org/wiki/Channing_Tatum
Charisma Carpenter	http://en.wikipedia.org/wiki/Charisma_Carpenter
Charlayne Hunter-Gault	http://en.wikipedia.org/wiki/Charlayne_Hunter-Gault
Charlemagne Palestine	http://en.wikipedia.org/wiki/Charlemagne_Palestine
Charlene Tilton	http://en.wikipedia.org/wiki/Charlene_Tilton
Charles "Buddy" Roemer III	http://en.wikipedia.org/wiki/Buddy_Roemer
Charles A. Graner	http://en.wikipedia.org/wiki/Charles_Graner
Charles A. Hayes	http://en.wikipedia.org/wiki/Charles_A._Hayes
Charles Abbott	http://en.wikipedia.org/wiki/Charles_Lydiard_Aubrey_Abbott
Charles Addams	http://en.wikipedia.org/wiki/Charles_Addams
Charles Augustin Sainte-Beuve	http://en.wikipedia.org/wiki/Charles_Augustin_Sainte-Beuve
Charles Aznavour	http://en.wikipedia.org/wiki/Charles_Aznavour
Charles B. Rangel	http://en.wikipedia.org/wiki/Charles_B._Rangel
Charles Babbage	http://en.wikipedia.org/wiki/Charles_Babbage
Charles Barkley	http://en.wikipedia.org/wiki/Charles_Barkley
Charles Batteux	http://en.wikipedia.org/wiki/Charles_Batteux
Charles Baudelaire	http://en.wikipedia.org/wiki/Charles_Baudelaire
Charles Bickford	http://en.wikipedia.org/wiki/Charles_Bickford
Charles Bonnet	http://en.wikipedia.org/wiki/Charles_Bonnet
Charles Boustany	http://en.wikipedia.org/wiki/Charles_Boustany
Charles Boyer	http://en.wikipedia.org/wiki/Charles_Boyer
Charles Boyle	http://en.wikipedia.org/wiki/Charles_Boyle,_4th_Earl_of_Orrery
Charles Bradlaugh	http://en.wikipedia.org/wiki/Charles_Bradlaugh
Charles Brockden Brown	http://en.wikipedia.org/wiki/Charles_Brockden_Brown
Charles Bronfman	http://en.wikipedia.org/wiki/Charles_Bronfman
Charles Bronson	http://en.wikipedia.org/wiki/Charles_Bronson
Charles Brown	http://en.wikipedia.org/wiki/Charles_Brown_(musician)
Charles Bukowski	http://en.wikipedia.org/wiki/Charles_Bukowski
Charles Bulfinch	http://en.wikipedia.org/wiki/Charles_Bulfinch
Charles Burney	http://en.wikipedia.org/wiki/Charles_Burney
Charles Burns	http://en.wikipedia.org/wiki/Charles_Burns_(cartoonist)
Charles C. Mann	http://en.wikipedia.org/wiki/Charles_C._Mann
Charles Canady	http://en.wikipedia.org/wiki/Charles_Canady
Charles Chesnutt	http://en.wikipedia.org/wiki/Charles_Chesnutt
Charles Churchill	http://en.wikipedia.org/wiki/Charles_Churchill_(satirist)
Charles Clarke	http://en.wikipedia.org/wiki/Charles_Clarke
Charles Coburn	http://en.wikipedia.org/wiki/Charles_Coburn
Charles Cornwallis	http://en.wikipedia.org/wiki/Charles_Cornwallis
Charles Cotesworth Pinckney	http://en.wikipedia.org/wiki/Charles_Cotesworth_Pinckney
Charles Cotton	http://en.wikipedia.org/wiki/Charles_Cotton
Charles Cullen	http://en.wikipedia.org/wiki/Charles_Cullen
Charles Curtis	http://en.wikipedia.org/wiki/Charles_Curtis
Charles Dance	http://en.wikipedia.org/wiki/Charles_Dance
Charles Darwin	http://en.wikipedia.org/wiki/Charles_Darwin
Charles de Gaulle	http://en.wikipedia.org/wiki/Charles_de_Gaulle
Charles de Lint	http://en.wikipedia.org/wiki/Charles_de_Lint
Charles Dibdin	http://en.wikipedia.org/wiki/Charles_Dibdin
Charles Dickens	http://en.wikipedia.org/wiki/Charles_Dickens
Charles Djou	http://en.wikipedia.org/wiki/Charles_Djou
Charles Drew	http://en.wikipedia.org/wiki/Charles_Drew
Charles Dudley Warner	http://en.wikipedia.org/wiki/Charles_Dudley_Warner
Charles Durning	http://en.wikipedia.org/wiki/Charles_Durning
Charles Dutton	http://en.wikipedia.org/wiki/Charles_S._Dutton
Charles E. Bennett	http://en.wikipedia.org/wiki/Charles_Edward_Bennett
Charles E. Merrill	http://en.wikipedia.org/wiki/Charles_E._Merrill
Charles E. Schumer	http://en.wikipedia.org/wiki/Charles_E._Schumer
Charles E. Whittaker	http://en.wikipedia.org/wiki/Charles_E._Whittaker
Charles E. Wilson	http://en.wikipedia.org/wiki/Charles_E._Wilson
Charles �douard Guillaume	http://en.wikipedia.org/wiki/Charles_%C3%89douard_Guillaume
Charles Edward Russell	http://en.wikipedia.org/wiki/Charles_Edward_Russell
Charles Eliot Norton	http://en.wikipedia.org/wiki/Charles_Eliot_Norton
Charles Elton	http://en.wikipedia.org/wiki/Charles_Sutherland_Elton
Charles Emory Smith	http://en.wikipedia.org/wiki/Charles_Emory_Smith
Charles Evans Hughes	http://en.wikipedia.org/wiki/Charles_Evans_Hughes
Charles F. Brannan	http://en.wikipedia.org/wiki/Charles_F._Brannan
Charles F. Brush	http://en.wikipedia.org/wiki/Charles_F._Brush
Charles F. Kettering	http://en.wikipedia.org/wiki/Charles_F._Kettering
Charles Ferguson Smith	http://en.wikipedia.org/wiki/Charles_Ferguson_Smith
Charles Follen Adams	http://en.wikipedia.org/wiki/Charles_Follen_Adams
Charles Fort	http://en.wikipedia.org/wiki/Charles_Fort
Charles Francis Adams	http://en.wikipedia.org/wiki/Charles_Francis_Adams,_Sr.
Charles Francis Adams, Jr.	http://en.wikipedia.org/wiki/Charles_Francis_Adams%2C_Jr.
Charles Fran�ois Dumouriez	http://en.wikipedia.org/wiki/Charles-Fran%C3%A7ois_Dumouriez
Charles Fran�ois Sturm	http://en.wikipedia.org/wiki/Charles_Fran%C3%A7ois_Sturm
Charles Fried	http://en.wikipedia.org/wiki/Charles_Fried
Charles G. Dawes	http://en.wikipedia.org/wiki/Charles_G._Dawes
Charles G. Koch	http://en.wikipedia.org/wiki/Charles_G._Koch
Charles G. Ross	http://en.wikipedia.org/wiki/Charles_N._Ross
Charles Gatewood	http://en.wikipedia.org/wiki/Charles_B._Gatewood
Charles Gibson	http://en.wikipedia.org/wiki/Charles_Gibson
Charles Gleyre	http://en.wikipedia.org/wiki/Charles_Gleyre
Charles Glover Barkla	http://en.wikipedia.org/wiki/Charles_Glover_Barkla
Charles Godfrey Leland	http://en.wikipedia.org/wiki/Charles_Godfrey_Leland
Charles Goodyear	http://en.wikipedia.org/wiki/Charles_Goodyear
Charles Gounod	http://en.wikipedia.org/wiki/Charles_Gounod
Charles Griffes	http://en.wikipedia.org/wiki/Charles_Griffes
Charles Grodin	http://en.wikipedia.org/wiki/Charles_Grodin
Charles Guiteau	http://en.wikipedia.org/wiki/Charles_Guiteau
Charles H. Bonesteel III	http://en.wikipedia.org/wiki/Charles_H._Bonesteel_III
Charles H. Percy	http://en.wikipedia.org/wiki/Charles_H._Percy
Charles H. Townes	http://en.wikipedia.org/wiki/Charles_H._Townes
Charles Haid	http://en.wikipedia.org/wiki/Charles_Haid
Charles Hatcher	http://en.wikipedia.org/wiki/Charles_Floyd_Hatcher
Charles Haughey	http://en.wikipedia.org/wiki/Charles_Haughey
Charles Hayward	http://en.wikipedia.org/wiki/Charles_Hayward
Charles Hendry	http://en.wikipedia.org/wiki/Charles_Hendry
Charles Horace Mayo	http://en.wikipedia.org/wiki/Charles_Horace_Mayo
Charles II	http://en.wikipedia.org/wiki/Charles_II_of_England
Charles III	http://en.wikipedia.org/wiki/Charles_III,_Prince_of_Monaco
Charles IV	http://en.wikipedia.org/wiki/Charles_IV_of_Spain
Charles Ives	http://en.wikipedia.org/wiki/Charles_Ives
Charles IX	http://en.wikipedia.org/wiki/Charles_IX_of_France
Charles J. Pedersen	http://en.wikipedia.org/wiki/Charles_J._Pedersen
Charles James Fox	http://en.wikipedia.org/wiki/Charles_James_Fox
Charles James Lever	http://en.wikipedia.org/wiki/Charles_James_Lever
Charles John Canning	http://en.wikipedia.org/wiki/Charles_John_Canning
Charles Keating	http://en.wikipedia.org/wiki/Charles_Keating
Charles Kennedy	http://en.wikipedia.org/wiki/Charles_Kennedy
Charles King	http://en.wikipedia.org/wiki/Charles_King_(actor)
Charles Konan Banny	http://en.wikipedia.org/wiki/Charles_Konan_Banny
Charles Krauthammer	http://en.wikipedia.org/wiki/Charles_Krauthammer
Charles Kuralt	http://en.wikipedia.org/wiki/Charles_Kuralt
Charles L. Terry, Jr.	http://en.wikipedia.org/wiki/Charles_L._Terry%2C_Jr.
Charles Lamb	http://en.wikipedia.org/wiki/Charles_Lamb_(writer)
Charles Lane	http://en.wikipedia.org/wiki/Charles_Lane_(actor)
Charles Laughton	http://en.wikipedia.org/wiki/Charles_Laughton
Charles Lindbergh	http://en.wikipedia.org/wiki/Charles_Lindbergh
Charles Lindbergh, Jr.	http://en.wikipedia.org/wiki/Charles_Lindbergh%2C_Jr.
Charles Lyell	http://en.wikipedia.org/wiki/Charles_Lyell
Charles M. Schwab	http://en.wikipedia.org/wiki/Charles_M._Schwab
Charles MacArthur	http://en.wikipedia.org/wiki/Charles_MacArthur
Charles Major	http://en.wikipedia.org/wiki/Charles_Major
Charles Manson	http://en.wikipedia.org/wiki/Charles_Manson
Charles Marriott	http://en.wikipedia.org/wiki/Charles_Marriott
Charles Martel	http://en.wikipedia.org/wiki/Charles_Martel
Charles Martin Smith	http://en.wikipedia.org/wiki/Charles_Martin_Smith
Charles Mathias	http://en.wikipedia.org/wiki/Charles_Mathias
Charles Mathias, Jr.	http://en.wikipedia.org/wiki/Charles_Mathias%2C_Jr.
Charles Maurice de Talleyrand	http://en.wikipedia.org/wiki/Charles_Maurice_de_Talleyrand
Charles McLean Andrews	http://en.wikipedia.org/wiki/Charles_McLean_Andrews
Charles Mingus	http://en.wikipedia.org/wiki/Charles_Mingus
Charles Moore	http://en.wikipedia.org/wiki/Charles_H._Moore
Charles Murray	http://en.wikipedia.org/wiki/Charles_Murray_(author)
Charles Nelson Reilly	http://en.wikipedia.org/wiki/Charles_Nelson_Reilly
Charles Ng	http://en.wikipedia.org/wiki/Charles_Ng
Charles O. Porter	http://en.wikipedia.org/wiki/Charles_O._Porter
Charles O. Prince	http://en.wikipedia.org/wiki/Charles_O._Prince
Charles Olson	http://en.wikipedia.org/wiki/Charles_Olson
Charles Osgood	http://en.wikipedia.org/wiki/Charles_Osgood
Charles Perrault	http://en.wikipedia.org/wiki/Charles_Perrault
Charles Pinckney	http://en.wikipedia.org/wiki/Charles_Pinckney_(governor)
Charles R. Jackson	http://en.wikipedia.org/wiki/Charles_R._Jackson
Charles R. Schwab	http://en.wikipedia.org/wiki/Charles_R._Schwab
Charles R. Walgreen	http://en.wikipedia.org/wiki/Charles_R._Walgreen
Charles Rangel	http://en.wikipedia.org/wiki/Charles_Rangel
Charles Rennie Mackintosh	http://en.wikipedia.org/wiki/Charles_Rennie_Mackintosh
Charles Rocket	http://en.wikipedia.org/wiki/Charles_Rocket
Charles Rosher	http://en.wikipedia.org/wiki/Charles_Rosher
Charles S. Johnson	http://en.wikipedia.org/wiki/Charles_S._Johnson
Charles Schulz	http://en.wikipedia.org/wiki/Charles_Schulz
Charles Schwab	http://en.wikipedia.org/wiki/Charles_R._Schwab
Charles Shaughnessy	http://en.wikipedia.org/wiki/Charles_Shaughnessy
Charles Simic	http://en.wikipedia.org/wiki/Charles_Simic
Charles Stanley	http://en.wikipedia.org/wiki/Charles_Stanley
Charles Starkweather	http://en.wikipedia.org/wiki/Charles_Starkweather
Charles Stewart Parnell	http://en.wikipedia.org/wiki/Charles_Stewart_Parnell
Charles Sturt	http://en.wikipedia.org/wiki/Charles_Sturt
Charles Sumner	http://en.wikipedia.org/wiki/Charles_Sumner
Charles Taylor	http://en.wikipedia.org/wiki/Charles_H._Taylor
Charles the Bald	http://en.wikipedia.org/wiki/Charles_the_Bald
Charles the Fat	http://en.wikipedia.org/wiki/Charles_the_Fat
Charles the Simple	http://en.wikipedia.org/wiki/Charles_the_Simple
Charles Thomas Newton	http://en.wikipedia.org/wiki/Charles_Thomas_Newton
Charles Thomson	http://en.wikipedia.org/wiki/Charles_Thomson
Charles Tupper	http://en.wikipedia.org/wiki/Charles_Tupper
Charles Turnbull	http://en.wikipedia.org/wiki/Charles_Turnbull
Charles V	http://en.wikipedia.org/wiki/Charles_V_of_France
Charles Van Doren	http://en.wikipedia.org/wiki/Charles_Van_Doren
Charles Vest	http://en.wikipedia.org/wiki/Charles_Vest
Charles VI	http://en.wikipedia.org/wiki/Charles_VI_of_France
Charles Vidor	http://en.wikipedia.org/wiki/Charles_Vidor
Charles VII	http://en.wikipedia.org/wiki/Charles_VII_of_France
Charles VIII	http://en.wikipedia.org/wiki/Charles_VIII_of_France
Charles W. Fairbanks	http://en.wikipedia.org/wiki/Charles_W._Fairbanks
Charles W. Freeman, Jr.	http://en.wikipedia.org/wiki/Charles_W._Freeman%2C_Jr.
Charles W. Socarides	http://en.wikipedia.org/wiki/Charles_W._Socarides
Charles W. Stenholm	http://en.wikipedia.org/wiki/Charles_W._Stenholm
Charles Walker	http://en.wikipedia.org/wiki/Charles_Walker_(British_politician)
Charles Walters	http://en.wikipedia.org/wiki/Charles_Walters
Charles Wheatstone	http://en.wikipedia.org/wiki/Charles_Wheatstone
Charles Whitley	http://en.wikipedia.org/wiki/Charles_Whitley
Charles Whitman	http://en.wikipedia.org/wiki/Charles_Whitman
Charles Willson Peale	http://en.wikipedia.org/wiki/Charles_Willson_Peale
Charles Wilson	http://en.wikipedia.org/wiki/Charles_Wilson_(Texas_politician)
Charles Wuorinen	http://en.wikipedia.org/wiki/Charles_Wuorinen
Charles X	http://en.wikipedia.org/wiki/Charles_X
Charles, Duke of Orl�ans	http://en.wikipedia.org/wiki/Charles%2C_duc_d%27Orl%C3%A9ans
Charles-Augustin de Coulomb	http://en.wikipedia.org/wiki/Charles-Augustin_de_Coulomb
Charles-Bernard Renouvier	http://en.wikipedia.org/wiki/Charles-Bernard_Renouvier
Charles-Fran�ois Daubigny	http://en.wikipedia.org/wiki/Charles-Fran%C3%A7ois_Daubigny
Charles-Marie Widor	http://en.wikipedia.org/wiki/Charles-Marie_Widor
Charley Pride	http://en.wikipedia.org/wiki/Charley_Pride
Charlie Bass	http://en.wikipedia.org/wiki/Charles_Bass
Charlie Bell	http://en.wikipedia.org/wiki/Charlie_Bell
Charlie Burchill	http://en.wikipedia.org/wiki/Charlie_Burchill
Charlie Byrd	http://en.wikipedia.org/wiki/Charlie_Byrd
Charlie Callas	http://en.wikipedia.org/wiki/Charlie_Callas
Charlie Chaplin	http://en.wikipedia.org/wiki/Charlie_Chaplin
Charlie Christian	http://en.wikipedia.org/wiki/Charlie_Christian
Charlie Daniels	http://en.wikipedia.org/wiki/Charlie_Daniels
Charlie Dent	http://en.wikipedia.org/wiki/Charlie_Dent
Charlie Elphicke	http://en.wikipedia.org/wiki/Charlie_Elphicke
Charlie Finley	http://en.wikipedia.org/wiki/Charlie_Finley
Charlie Gonzalez	http://en.wikipedia.org/wiki/Charlie_Gonzalez
Charlie Haden	http://en.wikipedia.org/wiki/Charlie_Haden
Charlie Hunnam	http://en.wikipedia.org/wiki/Charlie_Hunnam
Charlie Hunter	http://en.wikipedia.org/wiki/Charlie_Hunter
Charlie Kaufman	http://en.wikipedia.org/wiki/Charlie_Kaufman
Charlie Melancon	http://en.wikipedia.org/wiki/Charlie_Melancon
Charlie Murphy	http://en.wikipedia.org/wiki/Charlie_Murphy
Charlie Norwood	http://en.wikipedia.org/wiki/Charlie_Norwood
Charlie Parker	http://en.wikipedia.org/wiki/Charlie_Parker
Charlie Rose	http://en.wikipedia.org/wiki/Charlie_Rose
Charlie Sheen	http://en.wikipedia.org/wiki/Charlie_Sheen
Charlie Stenholm	http://en.wikipedia.org/wiki/Charlie_Stenholm
Charlie Trotter	http://en.wikipedia.org/wiki/Charlie_Trotter
Charlie Watts	http://en.wikipedia.org/wiki/Charlie_Watts
Charlie Wilson	http://en.wikipedia.org/wiki/Charlie_Wilson_(Ohio_politician)
Charlize Theron	http://en.wikipedia.org/wiki/Charlize_Theron
Charlotte Bront�	http://en.wikipedia.org/wiki/Charlotte_Bront%C3%AB
Charlotte Caffey	http://en.wikipedia.org/wiki/Charlotte_Caffey
Charlotte Church	http://en.wikipedia.org/wiki/Charlotte_Church
Charlotte Froom	http://en.wikipedia.org/wiki/Charlotte_Froom
Charlotte Leslie	http://en.wikipedia.org/wiki/Charlotte_Leslie
Charlotte MacLeod	http://en.wikipedia.org/wiki/Charlotte_MacLeod
Charlotte Perkins Gilman	http://en.wikipedia.org/wiki/Charlotte_Perkins_Gilman
Charlotte Rae	http://en.wikipedia.org/wiki/Charlotte_Rae
Charlotte Rampling	http://en.wikipedia.org/wiki/Charlotte_Rampling
Charlotte Ross	http://en.wikipedia.org/wiki/Charlotte_Ross
Charlotte von Stein	http://en.wikipedia.org/wiki/Charlotte_von_Stein
Charlton Heston	http://en.wikipedia.org/wiki/Charlton_Heston
Chastity Bono	http://en.wikipedia.org/wiki/Chastity_Bono
Chava Alberstein	http://en.wikipedia.org/wiki/Chava_Alberstein
Chazz Palminteri	http://en.wikipedia.org/wiki/Chazz_Palminteri
Che Guevara	http://en.wikipedia.org/wiki/Che_Guevara
Cheech Marin	http://en.wikipedia.org/wiki/Cheech_Marin
Chellie Pingree	http://en.wikipedia.org/wiki/Chellie_Pingree
Chelsea Clinton	http://en.wikipedia.org/wiki/Chelsea_Clinton
Chelsea Noble	http://en.wikipedia.org/wiki/Chelsea_Noble
Chely Wright	http://en.wikipedia.org/wiki/Chely_Wright
Chen Kenichi	http://en.wikipedia.org/wiki/Chen_Kenichi
Chen Ning Yang	http://en.wikipedia.org/wiki/Chen_Ning_Yang
Chen Shui-bian	http://en.wikipedia.org/wiki/Chen_Shui-bian
Cheri Oteri	http://en.wikipedia.org/wiki/Cheri_Oteri
Cherry Jones	http://en.wikipedia.org/wiki/Cherry_Jones
Cheryl Gillan	http://en.wikipedia.org/wiki/Cheryl_Gillan
Cheryl Hines	http://en.wikipedia.org/wiki/Cheryl_Hines
Cheryl Ladd	http://en.wikipedia.org/wiki/Cheryl_Ladd
Cheryl Lynn	http://en.wikipedia.org/wiki/Cheryl_Lynn
Cheryl Tiegs	http://en.wikipedia.org/wiki/Cheryl_Tiegs
Chesney Allen	http://en.wikipedia.org/wiki/Chesney_Allen
Chester A. Arthur	http://en.wikipedia.org/wiki/Chester_A._Arthur
Chester Bennington	http://en.wikipedia.org/wiki/Chester_Bennington
Chester Bowles	http://en.wikipedia.org/wiki/Chester_Bowles
Chester Brown	http://en.wikipedia.org/wiki/Chester_Brown
Chester G. Atkins	http://en.wikipedia.org/wiki/Chester_G._Atkins
Chester Gould	http://en.wikipedia.org/wiki/Chester_Gould
Chester Himes	http://en.wikipedia.org/wiki/Chester_Himes
Chester Kallman	http://en.wikipedia.org/wiki/Chester_Kallman
Chester W. Nimitz	http://en.wikipedia.org/wiki/Chester_W._Nimitz
Chet Allen	http://en.wikipedia.org/wiki/Chet_Allen
Chet Atkins	http://en.wikipedia.org/wiki/Chet_Atkins
Chet Baker	http://en.wikipedia.org/wiki/Chet_Baker
Chet Edwards	http://en.wikipedia.org/wiki/Chet_Edwards
Chet Huntley	http://en.wikipedia.org/wiki/Chet_Huntley
Chevy Chase	http://en.wikipedia.org/wiki/Chevy_Chase
Chi Chi La Rue	http://en.wikipedia.org/wiki/Chi_Chi_La_Rue
Chi Chi Rodriguez	http://en.wikipedia.org/wiki/Chi_Chi_Rodriguez
Chi McBride	http://en.wikipedia.org/wiki/Chi_McBride
Chiang Ching-Kuo	http://en.wikipedia.org/wiki/Chiang_Ching-Kuo
Chiang Kai-Shek	http://en.wikipedia.org/wiki/Chiang_Kai-Shek
Chic Hecht	http://en.wikipedia.org/wiki/Chic_Hecht
Chick Corea	http://en.wikipedia.org/wiki/Chick_Corea
Chico Marx	http://en.wikipedia.org/wiki/Chico_Marx
Chill Wills	http://en.wikipedia.org/wiki/Chill_Wills
Chino Moreno	http://en.wikipedia.org/wiki/Chino_Moreno
Chinua Achebe	http://en.wikipedia.org/wiki/Chinua_Achebe
Chinyelu Onwurah	http://en.wikipedia.org/wiki/Chinyelu_Onwurah
Chip E	http://en.wikipedia.org/wiki/Chip_E
Chip Kidd	http://en.wikipedia.org/wiki/Chip_Kidd
Chip Pashayan	http://en.wikipedia.org/wiki/Chip_Pashayan
Chip Pickering	http://en.wikipedia.org/wiki/Chip_Pickering
Chipper Jones	http://en.wikipedia.org/wiki/Chipper_Jones
Chirstopher Murphy	http://en.wikipedia.org/wiki/Christopher_murphy
Chita Rivera	http://en.wikipedia.org/wiki/Chita_Rivera
Chlodwig zu Hohenlohe-Schillingsfurst	http://en.wikipedia.org/wiki/Chlodwig_zu_Hohenlohe-Schillingsfurst
Chloe Sevigny	http://en.wikipedia.org/wiki/Chloe_Sevigny
Chloe Smith	http://en.wikipedia.org/wiki/Chloe_Smith
Choe Yong-rim	http://en.wikipedia.org/wiki/Choe_Yong-rim
Chopper Read	http://en.wikipedia.org/wiki/Chopper_Read
Choummaly Sayasone	http://en.wikipedia.org/wiki/Choummaly_Sayasone
Chow Yun-Fat	http://en.wikipedia.org/wiki/Chow_Yun-Fat
Chr�tien de Troyes	http://en.wikipedia.org/wiki/Chr%C3%A9tien_de_Troyes
Chris Alberghini	http://en.wikipedia.org/wiki/Chris_Alberghini
Chris Albers	http://en.wikipedia.org/wiki/Christijan_Albers
Chris Allen	http://en.wikipedia.org/wiki/Chris_Allen_%28footballer_born_1989%29
Chris Barrie	http://en.wikipedia.org/wiki/Chris_Barrie
Chris Bell	http://en.wikipedia.org/wiki/Chris_Bell_(politician)
Chris Botti	http://en.wikipedia.org/wiki/Chris_Botti
Chris Bryant	http://en.wikipedia.org/wiki/Chris_Bryant
Chris Burke	http://en.wikipedia.org/wiki/Chris_Burke_(actor)
Chris Cannon	http://en.wikipedia.org/wiki/Chris_Cannon
Chris Carmack	http://en.wikipedia.org/wiki/Chris_Carmack
Chris Carney	http://en.wikipedia.org/wiki/Chris_Carney
Chris Carter	http://en.wikipedia.org/wiki/Chris_Carter_%28left-handed_hitter%29
Chris Chocola	http://en.wikipedia.org/wiki/Chris_Chocola
Chris Columbus	http://en.wikipedia.org/wiki/Chris_Columbus_(filmmaker)
Chris Cooper	http://en.wikipedia.org/wiki/Chris_Cooper_(actor)
Chris Cornell	http://en.wikipedia.org/wiki/Chris_Cornell
Chris Cutler	http://en.wikipedia.org/wiki/Chris_Cutler
Chris Dodd	http://en.wikipedia.org/wiki/Chris_Dodd
Chris Elliott	http://en.wikipedia.org/wiki/Chris_Elliott
Chris Evans	http://en.wikipedia.org/wiki/Chris_Evans_(UK_politician)
Chris Evert	http://en.wikipedia.org/wiki/Chris_Evert
Chris Farley	http://en.wikipedia.org/wiki/Chris_Farley
Chris Frantz	http://en.wikipedia.org/wiki/Chris_Frantz
Chris Goss	http://en.wikipedia.org/wiki/Chris_Goss
Chris Grayling	http://en.wikipedia.org/wiki/Chris_Grayling
Chris Gregoire	http://en.wikipedia.org/wiki/Chris_Gregoire
Chris Heaton-Harris	http://en.wikipedia.org/wiki/Chris_Heaton-Harris
Chris Huhne	http://en.wikipedia.org/wiki/Chris_Huhne
Chris Isaak	http://en.wikipedia.org/wiki/Chris_Isaak
Chris Jeffs	http://en.wikipedia.org/wiki/Chris_Jeffs
Chris John	http://en.wikipedia.org/wiki/Chris_John
Chris Kattan	http://en.wikipedia.org/wiki/Chris_Kattan
Chris Kelly	http://en.wikipedia.org/wiki/Chris_Kelly_(British_politician)
Chris Kirkpatrick	http://en.wikipedia.org/wiki/Chris_Kirkpatrick
Chris Klein	http://en.wikipedia.org/wiki/Chris_Klein_(actor)
Chris Lambert	http://en.wikipedia.org/wiki/Chris_Lambert_(athlete)
Chris Langton	http://en.wikipedia.org/wiki/Chris_Langton
Chris Lee	http://en.wikipedia.org/wiki/Chris_Lee_(politician)
Chris Lowe	http://en.wikipedia.org/wiki/Chris_Lowe
Chris Makepeace	http://en.wikipedia.org/wiki/Chris_Makepeace
Chris Martin	http://en.wikipedia.org/wiki/Chris_Martin
Chris Masterson	http://en.wikipedia.org/wiki/Chris_Masterson
Chris Matthews	http://en.wikipedia.org/wiki/Chris_Matthews
Chris Moneymaker	http://en.wikipedia.org/wiki/Chris_Moneymaker
Chris Morris	http://en.wikipedia.org/wiki/Chris_Morris_(satirist)
Chris Noth	http://en.wikipedia.org/wiki/Chris_Noth
Chris O'Donnell	http://en.wikipedia.org/wiki/Chris_O%27Donnell
Chris Onstad	http://en.wikipedia.org/wiki/Chris_Onstad
Chris Parnell	http://en.wikipedia.org/wiki/Chris_Parnell
Chris Patten	http://en.wikipedia.org/wiki/Chris_Patten
Chris Pedersen	http://en.wikipedia.org/wiki/Chris_Pedersen_(musician)
Chris Penn	http://en.wikipedia.org/wiki/Chris_Penn
Chris Pine	http://en.wikipedia.org/wiki/Chris_Pine
Chris Pontius	http://en.wikipedia.org/wiki/Chris_Pontius
Chris Potter	http://en.wikipedia.org/wiki/Chris_Potter_(actor)
Chris Robinson	http://en.wikipedia.org/wiki/Chris_Robinson_(singer)
Chris Rock	http://en.wikipedia.org/wiki/Chris_Rock
Chris Ruane	http://en.wikipedia.org/wiki/Chris_Ruane
Chris Sarandon	http://en.wikipedia.org/wiki/Chris_Sarandon
Chris Skidmore	http://en.wikipedia.org/wiki/Chris_Skidmore
Chris Smith	http://en.wikipedia.org/wiki/Chris_Smith_(New_Jersey_politician)
Chris Squire	http://en.wikipedia.org/wiki/Chris_Squire
Chris Titus	http://en.wikipedia.org/wiki/Chris_Titus
Chris Tucker	http://en.wikipedia.org/wiki/Chris_Tucker
Chris van Abkoude	http://en.wikipedia.org/wiki/Chris_van_Abkoude
Chris Van Hollen	http://en.wikipedia.org/wiki/Chris_Van_Hollen
Chris Vrenna	http://en.wikipedia.org/wiki/Chris_Vrenna
Chris Wallace	http://en.wikipedia.org/wiki/Chris_Wallace_(journalist)
Chris Ware	http://en.wikipedia.org/wiki/Chris_Ware
Chris Watson	http://en.wikipedia.org/wiki/Chris_Watson
Chris Webber	http://en.wikipedia.org/wiki/Chris_Webber
Chris White	http://en.wikipedia.org/wiki/Chris_White_(politician)
Chris Whittle	http://en.wikipedia.org/wiki/Chris_Whittle
Chris Williamson	http://en.wikipedia.org/wiki/Chris_Williamson_(politician)
Chrissie Hynde	http://en.wikipedia.org/wiki/Chrissie_Hynde
Christa McAuliffe	http://en.wikipedia.org/wiki/Christa_McAuliffe
Christa Miller	http://en.wikipedia.org/wiki/Christa_Miller
Christa Wolf	http://en.wikipedia.org/wiki/Christa_Wolf
Christiaan Barnard	http://en.wikipedia.org/wiki/Christiaan_Barnard
Christiaan Huygens	http://en.wikipedia.org/wiki/Christiaan_Huygens
Christian Abt	http://en.wikipedia.org/wiki/Christian_Abt
Christian Alvart	http://en.wikipedia.org/wiki/Christian_Alvart
Christian Anfinsen	http://en.wikipedia.org/wiki/Christian_Anfinsen
Christian Bale	http://en.wikipedia.org/wiki/Christian_Bale
Christian Brando	http://en.wikipedia.org/wiki/Christian_Brando
Christian Campbell	http://en.wikipedia.org/wiki/Christian_Campbell
Christian Dior	http://en.wikipedia.org/wiki/Christian_Dior
Christian Doppler	http://en.wikipedia.org/wiki/Christian_Doppler
Christian Duguay	http://en.wikipedia.org/wiki/Christian_Duguay
Christian Herter	http://en.wikipedia.org/wiki/Christian_Herter
Christian Lacroix	http://en.wikipedia.org/wiki/Christian_Lacroix
Christian Lange	http://en.wikipedia.org/wiki/Christian_Lange
Christian Schwarz-Schilling	http://en.wikipedia.org/wiki/Christian_Schwarz-Schilling
Christian Slater	http://en.wikipedia.org/wiki/Christian_Slater
Christian Wolff	http://en.wikipedia.org/wiki/Christian_Wolff_(composer)
Christiane Amanpour	http://en.wikipedia.org/wiki/Christiane_Amanpour
Christie Brinkley	http://en.wikipedia.org/wiki/Christie_Brinkley
Christie Hefner	http://en.wikipedia.org/wiki/Christie_Hefner
Christina Aguilera	http://en.wikipedia.org/wiki/Christina_Aguilera
Christina Alessi	http://en.wikipedia.org/wiki/Christina_Alessi
Christina Applegate	http://en.wikipedia.org/wiki/Christina_Applegate
Christina Hoff Sommers	http://en.wikipedia.org/wiki/Christina_Hoff_Sommers
Christina Milian	http://en.wikipedia.org/wiki/Christina_Milian
Christina of Sweden	http://en.wikipedia.org/wiki/Christina_of_Sweden
Christina Onassis	http://en.wikipedia.org/wiki/Christina_Onassis
Christina Ricci	http://en.wikipedia.org/wiki/Christina_Ricci
Christina Rossetti	http://en.wikipedia.org/wiki/Christina_Rossetti
Christina Stead	http://en.wikipedia.org/wiki/Christina_Stead
Christine Baranski	http://en.wikipedia.org/wiki/Christine_Baranski
Christine Brooke-Rose	http://en.wikipedia.org/wiki/Christine_Brooke-Rose
Christine de Pizan	http://en.wikipedia.org/wiki/Christine_de_Pizan
Christine Elise	http://en.wikipedia.org/wiki/Christine_Elise
Christine Gregoire	http://en.wikipedia.org/wiki/Christine_Gregoire
Christine Jorgensen	http://en.wikipedia.org/wiki/Christine_Jorgensen
Christine Keeler	http://en.wikipedia.org/wiki/Christine_Keeler
Christine Lahti	http://en.wikipedia.org/wiki/Christine_Lahti
Christine Lakin	http://en.wikipedia.org/wiki/Christine_Lakin
Christine McVie	http://en.wikipedia.org/wiki/Christine_McVie
Christine Taylor	http://en.wikipedia.org/wiki/Christine_Taylor
Christine Todd Whitman	http://en.wikipedia.org/wiki/Christine_Todd_Whitman
Christoph Willibald Gluck	http://en.wikipedia.org/wiki/Christoph_Willibald_Gluck
Christopher Alexander	http://en.wikipedia.org/wiki/Christopher_Alexander
Christopher Atkins	http://en.wikipedia.org/wiki/Christopher_Atkins
Christopher Buckley	http://en.wikipedia.org/wiki/Christopher_Buckley
Christopher Chope	http://en.wikipedia.org/wiki/Christopher_Chope
Christopher Columbus	http://en.wikipedia.org/wiki/Christopher_Columbus
Christopher Cox	http://en.wikipedia.org/wiki/Christopher_Cox
Christopher Cross	http://en.wikipedia.org/wiki/Christopher_Cross
Christopher Eccleston	http://en.wikipedia.org/wiki/Christopher_Eccleston
Christopher George	http://en.wikipedia.org/wiki/Christopher_George
Christopher Guest	http://en.wikipedia.org/wiki/Christopher_Guest
Christopher H. Smith	http://en.wikipedia.org/wiki/Christopher_H._Smith
Christopher Hansteen	http://en.wikipedia.org/wiki/Christopher_Hansteen
Christopher Hewett	http://en.wikipedia.org/wiki/Christopher_Hewett
Christopher Hitchens	http://en.wikipedia.org/wiki/Christopher_Hitchens
Christopher Isherwood	http://en.wikipedia.org/wiki/Christopher_Isherwood
Christopher J. Dodd	http://en.wikipedia.org/wiki/Christopher_J._Dodd
Christopher Jones	http://en.wikipedia.org/wiki/Christopher_Jones_(actor)
Christopher Judge	http://en.wikipedia.org/wiki/Christopher_Judge
Christopher Knight	http://en.wikipedia.org/wiki/Christopher_Knight
Christopher Lambert	http://en.wikipedia.org/wiki/Christopher_Lambert
Christopher Lasch	http://en.wikipedia.org/wiki/Christopher_Lasch
Christopher Lee	http://en.wikipedia.org/wiki/Christopher_Lee
Christopher Leslie	http://en.wikipedia.org/wiki/Christopher_Leslie
Christopher Lloyd	http://en.wikipedia.org/wiki/Christopher_Lloyd
Christopher Lowell	http://en.wikipedia.org/wiki/Christopher_Lowell
Christopher Marlowe	http://en.wikipedia.org/wiki/Christopher_Marlowe
Christopher Meloni	http://en.wikipedia.org/wiki/Christopher_Meloni
Christopher Morley	http://en.wikipedia.org/wiki/Christopher_Morley
Christopher Pike	http://en.wikipedia.org/wiki/Christopher_Pike_(author)
Christopher Plummer	http://en.wikipedia.org/wiki/Christopher_Plummer
Christopher Reeve	http://en.wikipedia.org/wiki/Christopher_Reeve
Christopher Rich	http://en.wikipedia.org/wiki/Christopher_Rich_(actor)
Christopher Scarver	http://en.wikipedia.org/wiki/Christopher_Scarver
Christopher Shays	http://en.wikipedia.org/wiki/Christopher_Shays
Christopher Stasheff	http://en.wikipedia.org/wiki/Christopher_Stasheff
Christopher Walken	http://en.wikipedia.org/wiki/Christopher_Walken
Christopher Wren	http://en.wikipedia.org/wiki/Christopher_Wren
Christy Carlson Romano	http://en.wikipedia.org/wiki/Christy_Carlson_Romano
Christy Mathewson	http://en.wikipedia.org/wiki/Christy_Mathewson
Christy Turlington	http://en.wikipedia.org/wiki/Christy_Turlington
Chubby Checker	http://en.wikipedia.org/wiki/Chubby_Checker
Chuck Barris	http://en.wikipedia.org/wiki/Chuck_Barris
Chuck Berry	http://en.wikipedia.org/wiki/Chuck_Berry
Chuck Colson	http://en.wikipedia.org/wiki/Chuck_Colson
Chuck Connors	http://en.wikipedia.org/wiki/Chuck_Connors
Chuck D	http://en.wikipedia.org/wiki/Chuck_D
Chuck Forsberg	http://en.wikipedia.org/wiki/Chuck_Forsberg
Chuck Geschke	http://en.wikipedia.org/wiki/Chuck_Geschke
Chuck Grassley	http://en.wikipedia.org/wiki/Chuck_Grassley
Chuck Hagel	http://en.wikipedia.org/wiki/Chuck_Hagel
Chuck Hansen	http://en.wikipedia.org/wiki/Chuck_Hansen
Chuck Hoberman	http://en.wikipedia.org/wiki/Chuck_Hoberman
Chuck Jones	http://en.wikipedia.org/wiki/Chuck_Jones
Chuck Mangione	http://en.wikipedia.org/wiki/Chuck_Mangione
Chuck Negron	http://en.wikipedia.org/wiki/Chuck_Negron
Chuck Norris	http://en.wikipedia.org/wiki/Chuck_Norris
Chuck Palahniuk	http://en.wikipedia.org/wiki/Chuck_Palahniuk
Chuck Robb	http://en.wikipedia.org/wiki/Chuck_Robb
Chuck Schuldiner	http://en.wikipedia.org/wiki/Chuck_Schuldiner
Chuck Schumer	http://en.wikipedia.org/wiki/Chuck_Schumer
Chuck Swindoll	http://en.wikipedia.org/wiki/Chuck_Swindoll
Chuck Woolery	http://en.wikipedia.org/wiki/Chuck_Woolery
Chuck Yeager	http://en.wikipedia.org/wiki/Chuck_Yeager
Chuck Zito	http://en.wikipedia.org/wiki/Chuck_Zito
Chuka Umunna	http://en.wikipedia.org/wiki/Chuka_Umunna
Chun Doo Hwan	http://en.wikipedia.org/wiki/Chun_Doo_Hwan
Chung Un-chan	http://en.wikipedia.org/wiki/Chung_Un-chan
Cicely Tyson	http://en.wikipedia.org/wiki/Cicely_Tyson
Cid Corman	http://en.wikipedia.org/wiki/Cid_Corman
Cillian Murphy	http://en.wikipedia.org/wiki/Cillian_Murphy
Cindy Ambuehl	http://en.wikipedia.org/wiki/Cindy_Ambuehl
Cindy Cohn	http://en.wikipedia.org/wiki/Cindy_Cohn
Cindy Crawford	http://en.wikipedia.org/wiki/Cindy_Crawford
Cindy Jackson	http://en.wikipedia.org/wiki/Cindy_Jackson
Cindy Sheehan	http://en.wikipedia.org/wiki/Cindy_Sheehan
Cindy Williams	http://en.wikipedia.org/wiki/Cindy_Williams
Ciro Rodriguez	http://en.wikipedia.org/wiki/Ciro_Rodriguez
Claes Oldenburg	http://en.wikipedia.org/wiki/Claes_Oldenburg
Claiborne Pell	http://en.wikipedia.org/wiki/Claiborne_Pell
Claire Bloom	http://en.wikipedia.org/wiki/Claire_Bloom
Claire Danes	http://en.wikipedia.org/wiki/Claire_Danes
Claire Forlani	http://en.wikipedia.org/wiki/Claire_Forlani
Claire McCaskill	http://en.wikipedia.org/wiki/Claire_McCaskill
Claire Perry	http://en.wikipedia.org/wiki/Claire_Perry
Claire Trevor	http://en.wikipedia.org/wiki/Claire_Trevor
Clancy Brown	http://en.wikipedia.org/wiki/Clancy_Brown
Clara Allen	http://en.wikipedia.org/wiki/Clara_Forsythe_Allen
Clara Barton	http://en.wikipedia.org/wiki/Clara_Barton
Clara Bow	http://en.wikipedia.org/wiki/Clara_Bow
Clara Petacci	http://en.wikipedia.org/wiki/Clara_Petacci
Clara Schumann	http://en.wikipedia.org/wiki/Clara_Schumann
Clare Boothe Luce	http://en.wikipedia.org/wiki/Clare_Boothe_Luce
Clarence "Du" Burns	http://en.wikipedia.org/wiki/Du_Burns
Clarence Allen	http://en.wikipedia.org/wiki/Clarence_Ray_Allen
Clarence Brown	http://en.wikipedia.org/wiki/Clarence_Brown
Clarence Clemons	http://en.wikipedia.org/wiki/Clarence_Clemons
Clarence Darrow	http://en.wikipedia.org/wiki/Clarence_Darrow
Clarence Day	http://en.wikipedia.org/wiki/Clarence_Day
Clarence E. Miller	http://en.wikipedia.org/wiki/Clarence_E._Miller
Clarence E. Mulford	http://en.wikipedia.org/wiki/Clarence_E._Mulford
Clarence Page	http://en.wikipedia.org/wiki/Clarence_Page
Clarence Thomas	http://en.wikipedia.org/wiki/Clarence_Thomas
Clarence Williams III	http://en.wikipedia.org/wiki/Clarence_Williams_III
Clark Ashton Smith	http://en.wikipedia.org/wiki/Clark_Ashton_Smith
Clark Clifford	http://en.wikipedia.org/wiki/Clark_Clifford
Clark Gable	http://en.wikipedia.org/wiki/Clark_Gable
Clark L. Hull	http://en.wikipedia.org/wiki/Clark_L._Hull
Clark T. Randt	http://en.wikipedia.org/wiki/Clark_T._Randt
Claud Cockburn	http://en.wikipedia.org/wiki/Claud_Cockburn
Claude Adrien Helv�tius	http://en.wikipedia.org/wiki/Claude-Adrien_Helv%C3%A9tius
Claude Akins	http://en.wikipedia.org/wiki/Claude_Akins
Claude Allen	http://en.wikipedia.org/wiki/Claude_Allen
Claude Bernard	http://en.wikipedia.org/wiki/Claude_Bernard
Claude Brown	http://en.wikipedia.org/wiki/Claude_Brown
Claude Cohen-Tannoudji	http://en.wikipedia.org/wiki/Claude_Cohen-Tannoudji
Claude Debussy	http://en.wikipedia.org/wiki/Claude_Debussy
Claude Jutra	http://en.wikipedia.org/wiki/Claude_Jutra
Claude L�vi-Strauss	http://en.wikipedia.org/wiki/Claude_L%C3%A9vi-Strauss
Claude McKay	http://en.wikipedia.org/wiki/Claude_McKay
Claude Monet	http://en.wikipedia.org/wiki/Claude_Monet
Claude Pepper	http://en.wikipedia.org/wiki/Claude_Pepper
Claude Rains	http://en.wikipedia.org/wiki/Claude_Rains
Claude Shannon	http://en.wikipedia.org/wiki/Claude_Shannon
Claude Simon	http://en.wikipedia.org/wiki/Claude_Simon
Claude-Louis Berthollet	http://en.wikipedia.org/wiki/Claude-Louis_Berthollet
Claudette Colbert	http://en.wikipedia.org/wiki/Claudette_Colbert
Claudia Black	http://en.wikipedia.org/wiki/Claudia_Black
Claudia Cardinale	http://en.wikipedia.org/wiki/Claudia_Cardinale
Claudia Christian	http://en.wikipedia.org/wiki/Claudia_Christian
Claudia Schiffer	http://en.wikipedia.org/wiki/Claudia_Schiffer
Claudine Longet	http://en.wikipedia.org/wiki/Claudine_Longet
Claudine Schneider	http://en.wikipedia.org/wiki/Claudine_Schneider
Cl�udio Hummes	http://en.wikipedia.org/wiki/Cl%C3%A1udio_Hummes
Claudio Monteverdi	http://en.wikipedia.org/wiki/Claudio_Monteverdi
Claudius II Gothicus	http://en.wikipedia.org/wiki/Claudius_II_Gothicus
Claus von Bulow	http://en.wikipedia.org/wiki/Claus_von_Bulow
Claus von Stauffenberg	http://en.wikipedia.org/wiki/Claus_von_Stauffenberg
Clay Aiken	http://en.wikipedia.org/wiki/Clay_Aiken
Clayton K. Yeutter	http://en.wikipedia.org/wiki/Clayton_K._Yeutter
Clayton M. Jones	http://en.wikipedia.org/wiki/Clayton_M._Jones
Clayton Moore	http://en.wikipedia.org/wiki/Clayton_Moore
Clea DuVall	http://en.wikipedia.org/wiki/Clea_DuVall
Cleanth Brooks	http://en.wikipedia.org/wiki/Cleanth_Brooks
Cleavon Little	http://en.wikipedia.org/wiki/Cleavon_Little
Clement Attlee	http://en.wikipedia.org/wiki/Clement_Attlee
Clement Clarke Moore	http://en.wikipedia.org/wiki/Clement_Clarke_Moore
Cleo Moore	http://en.wikipedia.org/wiki/Cleo_Moore
Cliff Burton	http://en.wikipedia.org/wiki/Cliff_Burton
Cliff Gorman	http://en.wikipedia.org/wiki/Cliff_Gorman
Cliff Martinez	http://en.wikipedia.org/wiki/Cliff_Martinez
Cliff Richard	http://en.wikipedia.org/wiki/Cliff_Richard
Cliff Robertson	http://en.wikipedia.org/wiki/Cliff_Robertson
Cliff Stearns	http://en.wikipedia.org/wiki/Cliff_Stearns
Cliff Stoll	http://en.wikipedia.org/wiki/Cliff_Stoll
Cliff Williams	http://en.wikipedia.org/wiki/Cliff_Williams
Clifford A. Pickover	http://en.wikipedia.org/wiki/Clifford_A._Pickover
Clifford D. Simak	http://en.wikipedia.org/wiki/Clifford_D._Simak
Clifford G. Shull	http://en.wikipedia.org/wiki/Clifford_G._Shull
Clifford Geertz	http://en.wikipedia.org/wiki/Clifford_Geertz
Clifford Hansen	http://en.wikipedia.org/wiki/Clifford_Hansen
Clifford Holland	http://en.wikipedia.org/wiki/Clifford_Holland
Clifford Irving	http://en.wikipedia.org/wiki/Clifford_Irving
Clifford K. Berryman	http://en.wikipedia.org/wiki/Clifford_K._Berryman
Clifford Odets	http://en.wikipedia.org/wiki/Clifford_K._Berryman
Clifford Olson	http://en.wikipedia.org/wiki/Clifford_Olson
Clifton Davis	http://en.wikipedia.org/wiki/Clifton_Davis
Clifton Webb	http://en.wikipedia.org/wiki/Clifton_Webb
Clint Black	http://en.wikipedia.org/wiki/Clint_Black
Clint Eastwood	http://en.wikipedia.org/wiki/Clint_Eastwood
Clint Howard	http://en.wikipedia.org/wiki/Clint_Eastwood
Clint Walker	http://en.wikipedia.org/wiki/Clint_Walker
Clinton Davisson	http://en.wikipedia.org/wiki/Clinton_Davisson
Clive Barker	http://en.wikipedia.org/wiki/Clive_Barker
Clive Betts	http://en.wikipedia.org/wiki/Clive_Betts
Clive Cussler	http://en.wikipedia.org/wiki/Clive_Cussler
Clive Efford	http://en.wikipedia.org/wiki/Clive_Efford
Clive Owen	http://en.wikipedia.org/wiki/Clive_Owen
Clive Swift	http://en.wikipedia.org/wiki/Clive_Swift
Cloris Leachman	http://en.wikipedia.org/wiki/Cloris_Leachman
Clyde Barrow	http://en.wikipedia.org/wiki/Clyde_Barrow
Clyde Harold Smith	http://en.wikipedia.org/wiki/Clyde_Harold_Smith
Clyde Tolson	http://en.wikipedia.org/wiki/Clyde_Tolson
Coco Chanel	http://en.wikipedia.org/wiki/Coco_Chanel
Cofer Black	http://en.wikipedia.org/wiki/Cofer_Black
Cokie Roberts	http://en.wikipedia.org/wiki/Cokie_Roberts
Col Needham	http://en.wikipedia.org/wiki/Col_Needham
Col. Robert Morgan	http://en.wikipedia.org/wiki/Robert_K._Morgan
Colbert King	http://en.wikipedia.org/wiki/Colbert_King
Cole Hauser	http://en.wikipedia.org/wiki/Cole_Hauser
Cole Porter	http://en.wikipedia.org/wiki/Cole_Porter
Cole Sprouse	http://en.wikipedia.org/wiki/Cole_Sprouse
Coleen Gray	http://en.wikipedia.org/wiki/Coleen_Gray
Coleman Hawkins	http://en.wikipedia.org/wiki/Coleman_Hawkins
Coleman Young	http://en.wikipedia.org/wiki/Coleman_Young
Colin Campbell	http://en.wikipedia.org/wiki/Colin_Campbell_%28ice_hockey%29
Colin Farrell	http://en.wikipedia.org/wiki/Colin_Farrell
Colin Ferguson	http://en.wikipedia.org/wiki/Colin_Ferguson_(convict)
Colin Firth	http://en.wikipedia.org/wiki/Colin_Firth
Colin Greenwood	http://en.wikipedia.org/wiki/Colin_Greenwood
Colin Hanks	http://en.wikipedia.org/wiki/Colin_Hanks
Colin Hay	http://en.wikipedia.org/wiki/Colin_Hay
Colin MacInnes	http://en.wikipedia.org/wiki/Colin_MacInnes
Colin Mochrie	http://en.wikipedia.org/wiki/Colin_Mochrie
Colin Powell	http://en.wikipedia.org/wiki/Colin_Powell
Colin Quinn	http://en.wikipedia.org/wiki/Colin_Quinn
Colleen Atwood	http://en.wikipedia.org/wiki/Colleen_Atwood
Colleen Dewhurst	http://en.wikipedia.org/wiki/Colleen_Dewhurst
Colleen Kollar-Kotelly	http://en.wikipedia.org/wiki/Colleen_Kollar-Kotelly
Colley Cibber	http://en.wikipedia.org/wiki/Colley_Cibber
Collin Peterson	http://en.wikipedia.org/wiki/Collin_Peterson
Collin Walcott	http://en.wikipedia.org/wiki/Collin_Walcott
Colm Meaney	http://en.wikipedia.org/wiki/Collin_Walcott
Colm O'Ciosoig	http://en.wikipedia.org/wiki/Colm_O%27Ciosoig
Colonel Sanders	http://en.wikipedia.org/wiki/Colonel_Sanders
Colonel Tom Parker	http://en.wikipedia.org/wiki/Colonel_Tom_Parker
Columba Bush	http://en.wikipedia.org/wiki/Columba_Bush
Compay Segundo	http://en.wikipedia.org/wiki/Compay_Segundo
Compton MacKenzie	http://en.wikipedia.org/wiki/Compton_MacKenzie
Comte de Lautr�amont	http://en.wikipedia.org/wiki/Comte_de_Lautr%C3%A9amont
Conan O'Brien	http://en.wikipedia.org/wiki/Conan_O%27Brien
Conchata Ferrell	http://en.wikipedia.org/wiki/Conchata_Ferrell
Condoleezza Rice	http://en.wikipedia.org/wiki/Condoleezza_Rice
Connie Chung	http://en.wikipedia.org/wiki/Connie_Chung
Connie Francis	http://en.wikipedia.org/wiki/Connie_Francis
Connie Mack	http://en.wikipedia.org/wiki/Connie_Mack_III
Connie Mack	http://en.wikipedia.org/wiki/Connie_Mack_IV
Connie Mack	http://en.wikipedia.org/wiki/Connie_Mack_(baseball)
Connie Mack IV	http://en.wikipedia.org/wiki/Connie_Mack_IV
Connie Morella	http://en.wikipedia.org/wiki/Connie_Morella
Connie Nielsen	http://en.wikipedia.org/wiki/Connie_Nielsen
Connie Sellecca	http://en.wikipedia.org/wiki/Connie_Sellecca
Connie Stevens	http://en.wikipedia.org/wiki/Connie_Stevens
Connie Willis	http://en.wikipedia.org/wiki/Connie_Willis
Conor Burns	http://en.wikipedia.org/wiki/Conor_Burns
Conor Murphy	http://en.wikipedia.org/wiki/Conor_Murphy
Conor Oberst	http://en.wikipedia.org/wiki/Conor_Oberst
Conrad Aiken	http://en.wikipedia.org/wiki/Conrad_Aiken
Conrad Bain	http://en.wikipedia.org/wiki/Conrad_Bain
Conrad Black	http://en.wikipedia.org/wiki/Conrad_Black
Conrad Burns	http://en.wikipedia.org/wiki/Conrad_Burns
Conrad Hilton	http://en.wikipedia.org/wiki/Conrad_Hilton
Conrad Pellicanus	http://en.wikipedia.org/wiki/Conrad_Pellicanus
Conrad Richter	http://en.wikipedia.org/wiki/Conrad_Richter
Conrad Veidt	http://en.wikipedia.org/wiki/Conrad_Veidt
Constance Bennett	http://en.wikipedia.org/wiki/Constance_Bennett
Constance Cummings	http://en.wikipedia.org/wiki/Constance_Cummings
Constance Marie	http://en.wikipedia.org/wiki/Constance_Marie
Constance Moore	http://en.wikipedia.org/wiki/Constance_Moore
Constantin Brancusi	http://en.wikipedia.org/wiki/Constantin_Brancusi
Constantine the Great	http://en.wikipedia.org/wiki/Constantine_the_Great
Constantius II	http://en.wikipedia.org/wiki/Constantius_II
Conway Twitty	http://en.wikipedia.org/wiki/Conway_Twitty
Cookie Gilchrist	http://en.wikipedia.org/wiki/Cookie_Gilchrist
Cool Papa Bell	http://en.wikipedia.org/wiki/Cool_Papa_Bell
Cooper Evans	http://en.wikipedia.org/wiki/Cooper_Evans
Coral Eugene Watts	http://en.wikipedia.org/wiki/Coral_Eugene_Watts
Corazon Aquino	http://en.wikipedia.org/wiki/Corazon_Aquino
Corbin Bernsen	http://en.wikipedia.org/wiki/Corbin_Bernsen
Cordell Hull	http://en.wikipedia.org/wiki/Cordell_Hull
Coretta Scott King	http://en.wikipedia.org/wiki/Coretta_Scott_King
Coretta Scott King	http://en.wikipedia.org/wiki/Coretta_Scott_King
Corey Feldman	http://en.wikipedia.org/wiki/Corey_Feldman
Corey Haim	http://en.wikipedia.org/wiki/Corey_Haim
Corey Hart	http://en.wikipedia.org/wiki/Corey_Hart_(singer)
Corey Sevier	http://en.wikipedia.org/wiki/Corey_Sevier
Corey Taylor	http://en.wikipedia.org/wiki/Corey_Taylor
Corin Nemec	http://en.wikipedia.org/wiki/Corin_Nemec
Corin Redgrave	http://en.wikipedia.org/wiki/Corin_Redgrave
Corinne Calvet	http://en.wikipedia.org/wiki/Corinne_Calvet
Corinne Claiborne "Lindy" Boggs	http://en.wikipedia.org/wiki/Lindy_Boggs
Cormac McCarthy	http://en.wikipedia.org/wiki/Cormac_McCarthy
Cornel West	http://en.wikipedia.org/wiki/Cornel_West
Cornel Wilde	http://en.wikipedia.org/wiki/Cornel_Wilde
Cornelius Agrippa	http://en.wikipedia.org/wiki/Cornelius_Agrippa
Cornelius Cardew	http://en.wikipedia.org/wiki/Cornelius_Cardew
Cornelius Felton	http://en.wikipedia.org/wiki/Cornelius_Conway_Felton
Cornelius Gallus	http://en.wikipedia.org/wiki/Cornelius_Gallus
Cornelius Jansen	http://en.wikipedia.org/wiki/Cornelius_Jansen
Cornelius Janssen	http://en.wikipedia.org/wiki/Cornelius_Janssen
Cornelius Nepos	http://en.wikipedia.org/wiki/Cornelius_Nepos
Cornelius Vanderbilt	http://en.wikipedia.org/wiki/Cornelius_Vanderbilt
Cornell Woolrich	http://en.wikipedia.org/wiki/Cornell_Woolrich
Corrine Brown	http://en.wikipedia.org/wiki/Corrine_Brown
Cory Doctorow	http://en.wikipedia.org/wiki/Cory_Doctorow
Cory Wells	http://en.wikipedia.org/wiki/Cory_Wells
Cosey Fanni Tutti	http://en.wikipedia.org/wiki/Cosey_Fanni_Tutti
Cosimo de Medici	http://en.wikipedia.org/wiki/Cosimo_de_Medici
Costas Caramanlis	http://en.wikipedia.org/wiki/Costas_Caramanlis
Costas Caramanlis	http://en.wikipedia.org/wiki/Costas_Caramanlis
Costas Mandylor	http://en.wikipedia.org/wiki/Costas_Mandylor
Cotton Mather	http://en.wikipedia.org/wiki/Costas_Mandylor
Count Basie	http://en.wikipedia.org/wiki/Count_Basie
Countee Cullen	http://en.wikipedia.org/wiki/Countee_Cullen
Countess Vaughn	http://en.wikipedia.org/wiki/Countess_Vaughn
Country Joe McDonald	http://en.wikipedia.org/wiki/Country_Joe_McDonald
Courteney Cox	http://en.wikipedia.org/wiki/Courteney_Cox
Courtney B. Vance	http://en.wikipedia.org/wiki/Courtney_B._Vance
Courtney Love	http://en.wikipedia.org/wiki/Courtney_Love
Courtney Taylor	http://en.wikipedia.org/wiki/Courtney_Taylor-Taylor
Courtney Thorne-Smith	http://en.wikipedia.org/wiki/Courtney_Thorne-Smith
Coventry Patmore	http://en.wikipedia.org/wiki/Coventry_Patmore
Cozy Powell	http://en.wikipedia.org/wiki/Cozy_Powell
Craig Armstrong	http://en.wikipedia.org/wiki/Craig_Armstrong_(composer)
Craig Benson	http://en.wikipedia.org/wiki/Craig_Benson
Craig Bierko	http://en.wikipedia.org/wiki/Craig_Bierko
Craig Charles	http://en.wikipedia.org/wiki/Craig_Charles
Craig Crawford	http://en.wikipedia.org/wiki/Craig_Crawford
Craig David	http://en.wikipedia.org/wiki/Craig_David
Craig Ferguson	http://en.wikipedia.org/wiki/Craig_Ferguson
Craig Johnston	http://en.wikipedia.org/wiki/Craig_Johnston
Craig Kilborn	http://en.wikipedia.org/wiki/Craig_Kilborn
Craig McCracken	http://en.wikipedia.org/wiki/Craig_McCracken
Craig Mundie	http://en.wikipedia.org/wiki/Craig_Mundie
Craig Neidorf	http://en.wikipedia.org/wiki/Craig_Neidorf
Craig Newmark	http://en.wikipedia.org/wiki/Craig_Newmark
Craig Parker	http://en.wikipedia.org/wiki/Craig_Parker
Craig R. Barrett	http://en.wikipedia.org/wiki/Craig_R._Barrett
Craig Sheffer	http://en.wikipedia.org/wiki/Craig_Sheffer
Craig Shergold	http://en.wikipedia.org/wiki/Craig_Shergold
Craig Stevens	http://en.wikipedia.org/wiki/Craig_Stevens_(actor)
Craig T. Nelson	http://en.wikipedia.org/wiki/Craig_T._Nelson
Craig Thomas	http://en.wikipedia.org/wiki/Craig_L._Thomas
Craig Whittaker	http://en.wikipedia.org/wiki/Craig_Whittaker
Crazy Cabbie	http://en.wikipedia.org/wiki/Crazy_Cabbie
Crazy Horse	http://en.wikipedia.org/wiki/Crazy_Horse
Cree Summer	http://en.wikipedia.org/wiki/Cree_Summer
Creflo Dollar	http://en.wikipedia.org/wiki/Creflo_Dollar
Cresson H. Kearny	http://en.wikipedia.org/wiki/Cresson_H._Kearny
Cris Kirkwood	http://en.wikipedia.org/wiki/Cris_Kirkwood
Crispin Blunt	http://en.wikipedia.org/wiki/Crispin_Blunt
Crispin Glover	http://en.wikipedia.org/wiki/Crispin_Glover
Crispus Attucks	http://en.wikipedia.org/wiki/Crispus_Attucks
Criss Angel	http://en.wikipedia.org/wiki/Criss_Angel
Cristian Vogel	http://en.wikipedia.org/wiki/Cristian_Vogel
Cristiano Ronaldo	http://en.wikipedia.org/wiki/Cristiano_Ronaldo
Cristina Fern�ndez de Kirchner	http://en.wikipedia.org/wiki/Cristina_Fern%C3%A1ndez_de_Kirchner
Cristina Peri Rossi	http://en.wikipedia.org/wiki/Cristina_Peri_Rossi
Cristina Saralegui	http://en.wikipedia.org/wiki/Cristina_Saralegui
Crist�bal de Castillejo	http://en.wikipedia.org/wiki/Crist%C3%B3bal_de_Castillejo
Cruz Bustamante	http://en.wikipedia.org/wiki/Cruz_Bustamante
Crystal Bernard	http://en.wikipedia.org/wiki/Crystal_Bernard
Crystal Gayle	http://en.wikipedia.org/wiki/Crystal_Gayle
Crystal Waters	http://en.wikipedia.org/wiki/Crystal_Waters
Cuauhtemoc Cardenas	http://en.wikipedia.org/wiki/Cuauhtemoc_Cardenas
Cuba Gooding, Jr.	http://en.wikipedia.org/wiki/Cuba_Gooding%2C_Jr.
Curly Howard	http://en.wikipedia.org/wiki/Curly_Howard
Curt Flood	http://en.wikipedia.org/wiki/Curt_Flood
Curt Gowdy	http://en.wikipedia.org/wiki/Curt_Gowdy
Curt Schilling	http://en.wikipedia.org/wiki/Curt_Schilling
Curt Weldon	http://en.wikipedia.org/wiki/Curt_Weldon
Curtis Hanson	http://en.wikipedia.org/wiki/Curtis_Hanson
Curtis LeMay	http://en.wikipedia.org/wiki/Curtis_LeMay
Curtis Mayfield	http://en.wikipedia.org/wiki/Curtis_Mayfield
Curtis Sliwa	http://en.wikipedia.org/wiki/Curtis_Sliwa
Cushman Kellogg Davis	http://en.wikipedia.org/wiki/Cushman_Kellogg_Davis
Cy Young	http://en.wikipedia.org/wiki/Cy_Young
Cybill Shepherd	http://en.wikipedia.org/wiki/Cybill_Shepherd
Cyd Charisse	http://en.wikipedia.org/wiki/Cyd_Charisse
Cyndi Lauper	http://en.wikipedia.org/wiki/Cyndi_Lauper
Cynthia Geary	http://en.wikipedia.org/wiki/Cynthia_Geary
Cynthia Lummis	http://en.wikipedia.org/wiki/Cynthia_Lummis
Cynthia Macdonald	http://en.wikipedia.org/wiki/Cynthia_Macdonald
Cynthia McFadden	http://en.wikipedia.org/wiki/Cynthia_McFadden
Cynthia McKinney	http://en.wikipedia.org/wiki/Cynthia_McKinney
Cynthia Nixon	http://en.wikipedia.org/wiki/Cynthia_Nixon
Cynthia Ozick	http://en.wikipedia.org/wiki/Cynthia_Ozick
Cynthia Rowley	http://en.wikipedia.org/wiki/Cynthia_Rowley
Cynthia Weil	http://en.wikipedia.org/wiki/Cynthia_Weil
Cyrano de Bergerac	http://en.wikipedia.org/wiki/Cyrano_de_Bergerac
Cyril Connolly	http://en.wikipedia.org/wiki/Cyril_Connolly
Cyril Lucaris	http://en.wikipedia.org/wiki/Cyril_Lucaris
Cyril Neville	http://en.wikipedia.org/wiki/Cyril_Neville
Cyrus McCormick	http://en.wikipedia.org/wiki/Cyrus_McCormick
Cyrus the Great	http://en.wikipedia.org/wiki/Cyrus_the_Great
Cyrus Vance	http://en.wikipedia.org/wiki/Cyrus_Vance
Cyrus W. Field	http://en.wikipedia.org/wiki/Cyrus_W._Field
Czeslaw Milosz	http://en.wikipedia.org/wiki/Czeslaw_Milosz
D. B. Cooper	http://en.wikipedia.org/wiki/D._B._Cooper
D. B. Sweeney	http://en.wikipedia.org/wiki/D._B._Sweeney
D. French Slaughter, Jr.	http://en.wikipedia.org/wiki/D._French_Slaughter%2C_Jr.
D. H. Lawrence	http://en.wikipedia.org/wiki/D._H._Lawrence
D. L. Hughley	http://en.wikipedia.org/wiki/D._L._Hughley
D. M. Jayaratne	http://en.wikipedia.org/wiki/D._M._Jayaratne
D. W. Griffith	http://en.wikipedia.org/wiki/D._W._Griffith
Da Brat	http://en.wikipedia.org/wiki/Da_Brat
Dabney Coleman	http://en.wikipedia.org/wiki/Dabney_Coleman
Dack Rambo	http://en.wikipedia.org/wiki/Dack_Rambo
Daddy Yankee	http://en.wikipedia.org/wiki/Daddy_Yankee
Daevid Allen	http://en.wikipedia.org/wiki/Daevid_Allen
Dafydd ap Gwilym	http://en.wikipedia.org/wiki/Dafydd_ap_Gwilym
Dag Hammarskjold	http://en.wikipedia.org/wiki/Dag_Hammarskjold
Dagmar Krause	http://en.wikipedia.org/wiki/Dagmar_Krause
Dagobert I	http://en.wikipedia.org/wiki/Dagobert_I
Dahir Riyale Kahin	http://en.wikipedia.org/wiki/Dahir_Riyale_Kahin
Dai Havard	http://en.wikipedia.org/wiki/Dai_Havard
Daisy Berkowitz	http://en.wikipedia.org/wiki/Daisy_Berkowitz
Daisy Fuentes	http://en.wikipedia.org/wiki/Daisy_Fuentes
Dakota Fanning	http://en.wikipedia.org/wiki/Dakota_Fanning
Dalai Lama	http://en.wikipedia.org/wiki/14th_Dalai_Lama
Dale Bumpers	http://en.wikipedia.org/wiki/Dale_Bumpers
Dale Bumpers	http://en.wikipedia.org/wiki/Dale_Bumpers
Dale Carnegie	http://en.wikipedia.org/wiki/Dale_Carnegie
Dale Chihuly	http://en.wikipedia.org/wiki/Dale_Chihuly
Dale E. Kildee	http://en.wikipedia.org/wiki/Dale_E._Kildee
Dale E. Wolf	http://en.wikipedia.org/wiki/Dale_E._Wolf
Dale Earnhardt	http://en.wikipedia.org/wiki/Dale_Earnhardt
Dale Earnhardt, Jr.	http://en.wikipedia.org/wiki/Dale_Earnhardt%2C_Jr.
Dale Evans	http://en.wikipedia.org/wiki/Dale_Evans
Dale Kildee	http://en.wikipedia.org/wiki/Dale_Kildee
Dale Messick	http://en.wikipedia.org/wiki/Dale_Messick
Dale Midkiff	http://en.wikipedia.org/wiki/Dale_Midkiff
Dale Robertson	http://en.wikipedia.org/wiki/Dale_Robertson
Dalia Grybauskaitė	http://en.wikipedia.org/wiki/Dalia_Grybauskait%C4%97
Dalton Trumbo	http://en.wikipedia.org/wiki/Dalton_Trumbo
Dame Darcy	http://en.wikipedia.org/wiki/Dame_Darcy
Dame Pearlette Louisy	http://en.wikipedia.org/wiki/Dame_Pearlette_Louisy
Dame Silvia Cartwright	http://en.wikipedia.org/wiki/Dame_Silvia_Cartwright
Damian Collins	http://en.wikipedia.org/wiki/Damian_Collins
Damian Green	http://en.wikipedia.org/wiki/Damian_Green
Damian Hinds	http://en.wikipedia.org/wiki/Damian_Hinds
Damian Lewis	http://en.wikipedia.org/wiki/Damian_Lewis
Damien Hirst	http://en.wikipedia.org/wiki/Damien_Hirst
Damien Rice	http://en.wikipedia.org/wiki/Damien_Rice
Damo Suzuki	http://en.wikipedia.org/wiki/Damo_Suzuki
Damon Albarn	http://en.wikipedia.org/wiki/Damon_Albarn
Damon Dash	http://en.wikipedia.org/wiki/Damon_Dash
Damon Gough	http://en.wikipedia.org/wiki/Damon_Gough
Damon Runyon	http://en.wikipedia.org/wiki/Damon_Runyon
Damon Wayans	http://en.wikipedia.org/wiki/Damon_Wayans
Dan Abrams	http://en.wikipedia.org/wiki/Dan_Abrams
Dan Aykroyd	http://en.wikipedia.org/wiki/Dan_Aykroyd
Dan Balz	http://en.wikipedia.org/wiki/Dan_Balz
Dan Bartlett	http://en.wikipedia.org/wiki/Dan_Bartlett
Dan Blocker	http://en.wikipedia.org/wiki/Dan_Blocker
Dan Boren	http://en.wikipedia.org/wiki/Dan_Boren
Dan Brown	http://en.wikipedia.org/wiki/Dan_Brown
Dan Burton	http://en.wikipedia.org/wiki/Dan_Burton
Dan Burton	http://en.wikipedia.org/wiki/Dan_Burton
Dan Butler	http://en.wikipedia.org/wiki/Dan_Butler
Dan Castellaneta	http://en.wikipedia.org/wiki/Dan_Butler
Dan Castellaneta	http://en.wikipedia.org/wiki/Dan_Castellaneta
Dan Cortese	http://en.wikipedia.org/wiki/Dan_Cortese
Dan Dailey	http://en.wikipedia.org/wiki/Dan_Dailey
Dan Daniel	http://en.wikipedia.org/wiki/Dan_Daniel_(politician)
Dan Duryea	http://en.wikipedia.org/wiki/Dan_Duryea
Dan Farmer	http://en.wikipedia.org/wiki/Dan_Farmer
Dan Fogelberg	http://en.wikipedia.org/wiki/Dan_Fogelberg
Dan Fouts	http://en.wikipedia.org/wiki/Dan_Fouts
Dan Frisa	http://en.wikipedia.org/wiki/Dan_Frisa
Dan Futterman	http://en.wikipedia.org/wiki/Dan_Futterman
Dan Glickman	http://en.wikipedia.org/wiki/Dan_Glickman
Dan Glickman	http://en.wikipedia.org/wiki/Dan_Glickman
Dan Haggerty	http://en.wikipedia.org/wiki/Dan_Haggerty
Dan Harris	http://en.wikipedia.org/wiki/Dan_Harris
Dan Hedaya	http://en.wikipedia.org/wiki/Dan_Hedaya
Dan Lauria	http://en.wikipedia.org/wiki/Dan_Lauria
Dan Lipinski	http://en.wikipedia.org/wiki/Dan_Lipinski
Dan Lungren	http://en.wikipedia.org/wiki/Dan_Lungren
Dan Lungren	http://en.wikipedia.org/wiki/Dan_Lungren
Dan Maffei	http://en.wikipedia.org/wiki/Dan_Maffei
Dan Marino	http://en.wikipedia.org/wiki/Dan_Marino
Dan Miller	http://en.wikipedia.org/wiki/Dan_Miller_(U.S._politician)
Dan Moldea	http://en.wikipedia.org/wiki/Dan_Moldea
Dan O'Herlihy	http://en.wikipedia.org/wiki/Dan_O%27Herlihy
Dan Peek	http://en.wikipedia.org/wiki/Dan_Peek
Dan Penn	http://en.wikipedia.org/wiki/Dan_Penn
Dan Pink	http://en.wikipedia.org/wiki/Dan_Pink
Dan Quayle	http://en.wikipedia.org/wiki/Dan_Quayle
Dan Rather	http://en.wikipedia.org/wiki/Dan_Rather
Dan Rogerson	http://en.wikipedia.org/wiki/Dan_Rogerson
Dan Rostenkowski	http://en.wikipedia.org/wiki/Dan_Rostenkowski
Dan Rostenkowski	http://en.wikipedia.org/wiki/Dan_Rostenkowski
Dan Rowan	http://en.wikipedia.org/wiki/Dan_Rowan
Dan Savage	http://en.wikipedia.org/wiki/Dan_Rowan
Dan Schaefer	http://en.wikipedia.org/wiki/Dan_Rowan
Dan Schaefer	http://en.wikipedia.org/wiki/Dan_Schaefer
Dan Simmons	http://en.wikipedia.org/wiki/Dan_Simmons
Dan Snyder	http://en.wikipedia.org/wiki/Daniel_Snyder
Dan the Automator	http://en.wikipedia.org/wiki/Dan_the_Automator
Dan White	http://en.wikipedia.org/wiki/Dan_White
Dana Altman	http://en.wikipedia.org/wiki/Dana_Altman
Dana Andrews	http://en.wikipedia.org/wiki/Dana_Andrews
Dana Ashbrook	http://en.wikipedia.org/wiki/Dana_Ashbrook
Dana Carvey	http://en.wikipedia.org/wiki/Dana_Carvey
Dana Delany	http://en.wikipedia.org/wiki/Dana_Delany
Dana Elcar	http://en.wikipedia.org/wiki/Dana_Elcar
Dana Hill	http://en.wikipedia.org/wiki/Dana_Hill
Dana Ivey	http://en.wikipedia.org/wiki/Dana_Ivey
Dana Milbank	http://en.wikipedia.org/wiki/Dana_Milbank
Dana Plato	http://en.wikipedia.org/wiki/Dana_Plato
Dana Priest	http://en.wikipedia.org/wiki/Dana_Priest
Dana Reeve	http://en.wikipedia.org/wiki/Dana_Reeve
Dana Rohrabacher	http://en.wikipedia.org/wiki/Dana_Rohrabacher
Dana Snyder	http://en.wikipedia.org/wiki/Dana_Snyder
Dane Clark	http://en.wikipedia.org/wiki/Dane_Clark
Dane Cook	http://en.wikipedia.org/wiki/Dane_Cook
Dani Filth	http://en.wikipedia.org/wiki/Dani_Filth
Danica McKellar	http://en.wikipedia.org/wiki/Danica_McKellar
Danica Patrick	http://en.wikipedia.org/wiki/Danica_Patrick
Daniel A. Mica	http://en.wikipedia.org/wiki/Daniel_A._Mica
Daniel Acon	http://en.wikipedia.org/wiki/Daniel_Acon
Daniel Akaka	http://en.wikipedia.org/wiki/Daniel_Akaka
Daniel Alfredson	http://en.wikipedia.org/wiki/Daniel_Alfredson
Daniel Auber	http://en.wikipedia.org/wiki/Daniel-Fran%C3%A7ois-Esprit_Auber
Daniel Auteuil	http://en.wikipedia.org/wiki/Daniel_Auteuil
Daniel Bacon	http://en.wikipedia.org/wiki/Daniel_Bacon
Daniel Baldwin	http://en.wikipedia.org/wiki/Daniel_Baldwin
Daniel Bell	http://en.wikipedia.org/wiki/Daniel_Bell
Daniel Berrigan	http://en.wikipedia.org/wiki/Daniel_Berrigan
Daniel Boone	http://en.wikipedia.org/wiki/Daniel_Boone
Daniel Boorstin	http://en.wikipedia.org/wiki/Daniel_Boorstin
Daniel Byles	http://en.wikipedia.org/wiki/Daniel_Byles
Daniel C. Dennett	http://en.wikipedia.org/wiki/Daniel_C._Dennett
Daniel C. Tsui	http://en.wikipedia.org/wiki/Daniel_C._Tsui
Daniel Clowes	http://en.wikipedia.org/wiki/Daniel_Clowes
Daniel Craig	http://en.wikipedia.org/wiki/Daniel_Craig
Daniel D. Tompkins	http://en.wikipedia.org/wiki/Daniel_D._Tompkins
Daniel Dae Kim	http://en.wikipedia.org/wiki/Daniel_Dae_Kim
Daniel Davis	http://en.wikipedia.org/wiki/Daniel_Davis
Daniel Day-Lewis	http://en.wikipedia.org/wiki/Daniel_Day-Lewis
Daniel Defoe	http://en.wikipedia.org/wiki/Daniel_Defoe
Daniel Ellsberg	http://en.wikipedia.org/wiki/Daniel_Ellsberg
Daniel Ernst Jablonski	http://en.wikipedia.org/wiki/Daniel_Ernst_Jablonski
Daniel Inouye	http://en.wikipedia.org/wiki/Daniel_Inouye
Daniel J. Bernstein	http://en.wikipedia.org/wiki/Daniel_J._Bernstein
Daniel J. Evans	http://en.wikipedia.org/wiki/Daniel_J._Evans
Daniel J. Travanti	http://en.wikipedia.org/wiki/Daniel_J._Travanti
Daniel Johns	http://en.wikipedia.org/wiki/Daniel_Johns
Daniel K. Akaka	http://en.wikipedia.org/wiki/Daniel_K._Akaka
Daniel K. Inouye	http://en.wikipedia.org/wiki/Daniel_K._Inouye
Daniel Kawczynski	http://en.wikipedia.org/wiki/Daniel_Kawczynski
Daniel Keys Moran	http://en.wikipedia.org/wiki/Daniel_Keys_Moran
Daniel Mann	http://en.wikipedia.org/wiki/Daniel_Mann
Daniel Massey	http://en.wikipedia.org/wiki/Daniel_Massey_(actor)
Daniel O'Connell	http://en.wikipedia.org/wiki/Daniel_O%27Connell
Daniel Ortega	http://en.wikipedia.org/wiki/Daniel_Ortega
Daniel Patrick Moynihan	http://en.wikipedia.org/wiki/Daniel_Patrick_Moynihan
Daniel Patrick Moynihan	http://en.wikipedia.org/wiki/Daniel_Patrick_Moynihan
Daniel Pearl	http://en.wikipedia.org/wiki/Daniel_Pearl
Daniel Petrie	http://en.wikipedia.org/wiki/Daniel_Petrie
Daniel Pinkwater	http://en.wikipedia.org/wiki/Daniel_Pinkwater
Daniel Pipes	http://en.wikipedia.org/wiki/Daniel_Pipes
Daniel Poulter	http://en.wikipedia.org/wiki/Daniel_Poulter
Daniel R. Coats	http://en.wikipedia.org/wiki/Daniel_R._Coats
Daniel Radcliffe	http://en.wikipedia.org/wiki/Daniel_Radcliffe
Daniel Schorr	http://en.wikipedia.org/wiki/Daniel_Schorr
Daniel Shays	http://en.wikipedia.org/wiki/Daniel_Shays
Daniel Smith	http://en.wikipedia.org/wiki/Daniel_Wayne_Smith
Daniel Stern	http://en.wikipedia.org/wiki/Daniel_Stern_(actor)
Daniel Vierge	http://en.wikipedia.org/wiki/Daniel_Vierge
Daniel W. Bell	http://en.wikipedia.org/wiki/Daniel_W._Bell
Daniel Webster	http://en.wikipedia.org/wiki/Daniel_Webster
Daniel Yergin	http://en.wikipedia.org/wiki/Daniel_Yergin
Daniela Hantuchova	http://en.wikipedia.org/wiki/Daniela_Hantuchova
Daniela Pestova	http://en.wikipedia.org/wiki/Daniela_Pestova
Daniele Gaither	http://en.wikipedia.org/wiki/Daniele_Gaither
Danielle Berry	http://en.wikipedia.org/wiki/Danielle_Berry
Danielle Darrieux	http://en.wikipedia.org/wiki/Danielle_Darrieux
Danielle Dax	http://en.wikipedia.org/wiki/Danielle_Dax
Danielle Fishel	http://en.wikipedia.org/wiki/Danielle_Fishel
Danielle Harris	http://en.wikipedia.org/wiki/Danielle_Harris
Danielle Panabaker	http://en.wikipedia.org/wiki/Danielle_Panabaker
Danielle Steel	http://en.wikipedia.org/wiki/Danielle_Steel
Danilo T�rk	http://en.wikipedia.org/wiki/Danilo_T%C3%BCrk
Daniyal Akhmetov	http://en.wikipedia.org/wiki/Daniyal_Akhmetov
Dann Florek	http://en.wikipedia.org/wiki/Dann_Florek
Dannie Abse	http://en.wikipedia.org/wiki/Dannie_Abse
Dannii Minogue	http://en.wikipedia.org/wiki/Dannii_Minogue
Danny Aiello	http://en.wikipedia.org/wiki/Danny_Aiello
Danny Alexander	http://en.wikipedia.org/wiki/Danny_Alexander
Danny Bonaduce	http://en.wikipedia.org/wiki/Danny_Bonaduce
Danny Boyle	http://en.wikipedia.org/wiki/Danny_Boyle
Danny Carey	http://en.wikipedia.org/wiki/Danny_Carey
Danny Collins	http://en.wikipedia.org/wiki/Danny_Collins
Danny Davis	http://en.wikipedia.org/wiki/Danny_K._Davis
Danny DeVito	http://en.wikipedia.org/wiki/Danny_DeVito
Danny Elfman	http://en.wikipedia.org/wiki/Danny_Elfman
Danny Glover	http://en.wikipedia.org/wiki/Danny_Glover
Danny Hutton	http://en.wikipedia.org/wiki/Danny_Hutton
Danny Joe Brown	http://en.wikipedia.org/wiki/Danny_Joe_Brown
Danny Kaye	http://en.wikipedia.org/wiki/Danny_Kaye
Danny Lohner	http://en.wikipedia.org/wiki/Danny_Lohner
Danny Masterson	http://en.wikipedia.org/wiki/Danny_Masterson
Danny Pintauro	http://en.wikipedia.org/wiki/Danny_Pintauro
Danny Sugerman	http://en.wikipedia.org/wiki/Danny_Sugerman
Danny Thomas	http://en.wikipedia.org/wiki/Danny_Thomas
Danny Trejo	http://en.wikipedia.org/wiki/Danny_Trejo
Dante B. Fascell	http://en.wikipedia.org/wiki/Dante_B._Fascell
Dante Fascell	http://en.wikipedia.org/wiki/Dante_Fascell
Dante Gabriel Rossetti	http://en.wikipedia.org/wiki/Dante_Gabriel_Rossetti
Dante Hall	http://en.wikipedia.org/wiki/Dante_Hall
Daphne Du Maurier	http://en.wikipedia.org/wiki/Daphne_Du_Maurier
Daphne Zuniga	http://en.wikipedia.org/wiki/Daphne_Zuniga
Darby Crash	http://en.wikipedia.org/wiki/Darby_Crash
Darcy LaPier	http://en.wikipedia.org/wiki/Darcy_LaPier
D'arcy Wretzky	http://en.wikipedia.org/wiki/D%27arcy_Wretzky
Dario Argento	http://en.wikipedia.org/wiki/Dario_Argento
Dario Fo	http://en.wikipedia.org/wiki/Dario_Fo
Darius II Ochus	http://en.wikipedia.org/wiki/Darius_II_Ochus
Darius III Codomannus	http://en.wikipedia.org/wiki/Darius_III_Codomannus
Darius Milhaud	http://en.wikipedia.org/wiki/Darius_Milhaud
Darius Rucker	http://en.wikipedia.org/wiki/Darius_Rucker
Darius the Great	http://en.wikipedia.org/wiki/Darius_the_Great
Darl McBride	http://en.wikipedia.org/wiki/Darl_McBride
Darla Hood	http://en.wikipedia.org/wiki/Darla_Hood
Darlene Cates	http://en.wikipedia.org/wiki/Darlene_Cates
Darlene Hooley	http://en.wikipedia.org/wiki/Darlene_Hooley
Darlie Routier	http://en.wikipedia.org/wiki/Darlie_Routier
Daron Malakian	http://en.wikipedia.org/wiki/Daron_Malakian
Darrell Hammond	http://en.wikipedia.org/wiki/Darrell_Hammond
Darrell Issa	http://en.wikipedia.org/wiki/Darrell_Issa
Darrell Johnson	http://en.wikipedia.org/wiki/Darrell_Johnson
Darren Aronofsky	http://en.wikipedia.org/wiki/Darren_Aronofsky
Darren E. Burrows	http://en.wikipedia.org/wiki/Darren_E._Burrows
Darren Emerson	http://en.wikipedia.org/wiki/Darren_Emerson
Darren Hayes	http://en.wikipedia.org/wiki/Darren_Hayes
Darren McGavin	http://en.wikipedia.org/wiki/Darren_McGavin
Darryl F. Zanuck	http://en.wikipedia.org/wiki/Darryl_F._Zanuck
Darryl Strawberry	http://en.wikipedia.org/wiki/Darryl_Strawberry
Darva Conger	http://en.wikipedia.org/wiki/Darva_Conger
Daryl Gates	http://en.wikipedia.org/wiki/Daryl_Gates
Daryl Hall	http://en.wikipedia.org/wiki/Daryl_Hall
Daryl Hannah	http://en.wikipedia.org/wiki/Daryl_Hannah
Daryn Kagan	http://en.wikipedia.org/wiki/Daryn_Kagan
Dashiell Hammett	http://en.wikipedia.org/wiki/Dashiell_Hammett
Dave Abbruzzese	http://en.wikipedia.org/wiki/Dave_Abbruzzese
Dave Allen	http://en.wikipedia.org/wiki/Dave_Allen_(actor)
Dave Attell	http://en.wikipedia.org/wiki/Dave_Attell
Dave Barry	http://en.wikipedia.org/wiki/Dave_Barry
Dave Batista	http://en.wikipedia.org/wiki/Dave_Batista
Dave Blood	http://en.wikipedia.org/wiki/Dave_Blood
Dave Brubeck	http://en.wikipedia.org/wiki/Dave_Brubeck
Dave Camp	http://en.wikipedia.org/wiki/Dave_Camp
Dave Chappelle	http://en.wikipedia.org/wiki/Dave_Chappelle
Dave Clark	http://en.wikipedia.org/wiki/Dave_Clark_(musician)
Dave Coulier	http://en.wikipedia.org/wiki/Dave_Coulier
Dave Coverly	http://en.wikipedia.org/wiki/Dave_Coverly
Dave Davies	http://en.wikipedia.org/wiki/Dave_Davies
Dave Durenberger	http://en.wikipedia.org/wiki/Dave_Durenberger
Dave Edmunds	http://en.wikipedia.org/wiki/Dave_Edmunds
Dave Eggers	http://en.wikipedia.org/wiki/Dave_Eggers
Dave Foley	http://en.wikipedia.org/wiki/Dave_Foley
Dave Freudenthal	http://en.wikipedia.org/wiki/Dave_Freudenthal
Dave Freudenthal	http://en.wikipedia.org/wiki/Dave_Freudenthal
Dave Gahan	http://en.wikipedia.org/wiki/Dave_Gahan
Dave Garroway	http://en.wikipedia.org/wiki/Dave_Garroway
Dave Goodman	http://en.wikipedia.org/wiki/Dave_Goodman
Dave Greenslade	http://en.wikipedia.org/wiki/Dave_Greenslade
Dave Grohl	http://en.wikipedia.org/wiki/Dave_Grohl
Dave Heineman	http://en.wikipedia.org/wiki/Dave_Heineman
Dave Heineman	http://en.wikipedia.org/wiki/Dave_Heineman
Dave Kopay	http://en.wikipedia.org/wiki/Dave_Kopay
Dave Lebling	http://en.wikipedia.org/wiki/Dave_Lebling
Dave Loebsack	http://en.wikipedia.org/wiki/Dave_Loebsack
Dave Lombardo	http://en.wikipedia.org/wiki/Dave_Lombardo
Dave Matthews	http://en.wikipedia.org/wiki/Dave_Matthews
Dave McCurdy	http://en.wikipedia.org/wiki/Dave_McCurdy
Dave Mustaine	http://en.wikipedia.org/wiki/Dave_Mustaine
Dave Navarro	http://en.wikipedia.org/wiki/Dave_Navarro
Dave Pirner	http://en.wikipedia.org/wiki/Dave_Pirner
Dave Reichert	http://en.wikipedia.org/wiki/Dave_Reichert
Dave Riley	http://en.wikipedia.org/wiki/Dave_Riley
Dave Rowntree	http://en.wikipedia.org/wiki/Dave_Rowntree
Dave Sim	http://en.wikipedia.org/wiki/Dave_Sim
Dave Stewart	http://en.wikipedia.org/wiki/Dave_Stewart_(keyboardist)
Dave Stewart	http://en.wikipedia.org/wiki/David_A._Stewart
Dave Thomas	http://en.wikipedia.org/wiki/Dave_Thomas_(American_businessman)
Dave Watts	http://en.wikipedia.org/wiki/David_Watts_(politician)
Dave Weldon	http://en.wikipedia.org/wiki/Dave_Weldon
Dave Willis	http://en.wikipedia.org/wiki/Dave_Willis
Dave Winer	http://en.wikipedia.org/wiki/Dave_Winer
Dave Winfield	http://en.wikipedia.org/wiki/Dave_Winfield
Davey Havok	http://en.wikipedia.org/wiki/Davey_Havok
David A. Paterson	http://en.wikipedia.org/wiki/David_A._Paterson
David Abshire	http://en.wikipedia.org/wiki/David_Abshire
David Acomba	http://en.wikipedia.org/wiki/David_Acomba
David Addington	http://en.wikipedia.org/wiki/David_Addington
David Alan Grier	http://en.wikipedia.org/wiki/David_Alan_Grier
David Allan Coe	http://en.wikipedia.org/wiki/David_Allan_Coe
David Amess	http://en.wikipedia.org/wiki/David_Amess
David Anderson	http://en.wikipedia.org/wiki/David_Anderson_(UK_politician)
David Antin	http://en.wikipedia.org/wiki/David_Antin
David Arquette	http://en.wikipedia.org/wiki/David_Arquette
David Attenborough	http://en.wikipedia.org/wiki/David_Attenborough
David Axelrod	http://en.wikipedia.org/wiki/David_Axelrod
David B. Rivkin	http://en.wikipedia.org/wiki/David_B._Rivkin
David Baldacci	http://en.wikipedia.org/wiki/David_Baldacci
David Baltimore	http://en.wikipedia.org/wiki/David_Baltimore
David Banner	http://en.wikipedia.org/wiki/David_Banner
David Barton	http://en.wikipedia.org/wiki/David_Barton
David Beaton	http://en.wikipedia.org/wiki/David_Barton
David Beaty	http://en.wikipedia.org/wiki/David_Beaty
David Beckham	http://en.wikipedia.org/wiki/David_Beckham
David Belasco	http://en.wikipedia.org/wiki/David_Belasco
David Benedictus	http://en.wikipedia.org/wiki/David_Benedictus
David Ben-Gurion	http://en.wikipedia.org/wiki/David_Ben-Gurion
David Berkowitz	http://en.wikipedia.org/wiki/David_Berkowitz
David Bisbal	http://en.wikipedia.org/wiki/David_Bisbal
David Blaine	http://en.wikipedia.org/wiki/David_Blaine
David Bloom	http://en.wikipedia.org/wiki/David_Bloom
David Blunkett	http://en.wikipedia.org/wiki/David_Blunkett
David Bohm	http://en.wikipedia.org/wiki/David_Bohm
David Boies	http://en.wikipedia.org/wiki/David_Boies
David Bonior	http://en.wikipedia.org/wiki/David_Bonior
David Boreanaz	http://en.wikipedia.org/wiki/David_Boreanaz
David Bowie	http://en.wikipedia.org/wiki/David_Bowie
David Brancaccio	http://en.wikipedia.org/wiki/David_Brancaccio
David Brenner	http://en.wikipedia.org/wiki/David_Brenner
David Brin	http://en.wikipedia.org/wiki/David_Brin
David Brinkley	http://en.wikipedia.org/wiki/David_Brinkley
David Brock	http://en.wikipedia.org/wiki/David_Brock
David Broder	http://en.wikipedia.org/wiki/David_Broder
David Brooks	http://en.wikipedia.org/wiki/David_Brooks_(journalist)
David Brudnoy	http://en.wikipedia.org/wiki/David_Brudnoy
David Burke	http://en.wikipedia.org/wiki/David_Burke_(actor)
David Burrowes	http://en.wikipedia.org/wiki/David_Burrowes
David Burtka	http://en.wikipedia.org/wiki/David_Burtka
David Butler	http://en.wikipedia.org/wiki/David_Butler_(director)
David Byrne	http://en.wikipedia.org/wiki/David_Byrne
David C. Novak	http://en.wikipedia.org/wiki/David_C._Novak
David Cairns	http://en.wikipedia.org/wiki/David_Cairns_(politician)
David Cameron	http://en.wikipedia.org/wiki/David_Cameron
David Cannadine	http://en.wikipedia.org/wiki/David_Cannadine
David Carradine	http://en.wikipedia.org/wiki/David_Carradine
David Caruso	http://en.wikipedia.org/wiki/David_Caruso
David Cassidy	http://en.wikipedia.org/wiki/David_Cassidy
David Chalmers	http://en.wikipedia.org/wiki/David_Chalmers
David Charvet	http://en.wikipedia.org/wiki/David_Charvet
David Chokachi	http://en.wikipedia.org/wiki/David_Chokachi
David Copperfield	http://en.wikipedia.org/wiki/David_Copperfield_(illusionist)
David Coverdale	http://en.wikipedia.org/wiki/David_Coverdale
David Crane	http://en.wikipedia.org/wiki/David_Crane_(writer/producer)
David Crausby	http://en.wikipedia.org/wiki/David_Crausby
David Cronenberg	http://en.wikipedia.org/wiki/David_Cronenberg
David Crosby	http://en.wikipedia.org/wiki/David_Crosby
David Cross	http://en.wikipedia.org/wiki/David_Cross
David Cunningham	http://en.wikipedia.org/wiki/David_Cunningham_(musician)
David D. Smith	http://en.wikipedia.org/wiki/David_D._Smith
David Davies	http://en.wikipedia.org/wiki/Dave_Davies_%28Ontario_politician%29
David Davis	http://en.wikipedia.org/wiki/David_Davis_(British_politician)
David Desrosiers	http://en.wikipedia.org/wiki/David_Desrosiers
David Dinkins	http://en.wikipedia.org/wiki/David_Dinkins
David Doyle	http://en.wikipedia.org/wiki/David_Doyle_(actor)
David Dreier	http://en.wikipedia.org/wiki/David_Dreier
David Dreier	http://en.wikipedia.org/wiki/David_Dreier
David Duchovny	http://en.wikipedia.org/wiki/David_Duchovny
David Dudley Field	http://en.wikipedia.org/wiki/David_Dudley_Field
David Duke	http://en.wikipedia.org/wiki/David_Duke
David Dukes	http://en.wikipedia.org/wiki/David_Dukes
David Durenberger	http://en.wikipedia.org/wiki/David_Durenberger
David E. Bonior	http://en.wikipedia.org/wiki/David_E._Bonior
David E. Kelley	http://en.wikipedia.org/wiki/David_E._Kelley
David Eddings	http://en.wikipedia.org/wiki/David_Eddings
David Edward Maust	http://en.wikipedia.org/wiki/David_Edward_Maust
David Einhorn	http://en.wikipedia.org/wiki/David_Einhorn_(rabbi)
David Evennett	http://en.wikipedia.org/wiki/David_Evennett
David Farragut	http://en.wikipedia.org/wiki/David_Farragut
David Faustino	http://en.wikipedia.org/wiki/David_Faustino
David Filo	http://en.wikipedia.org/wiki/David_Filo
David Fincher	http://en.wikipedia.org/wiki/David_Fincher
David Foster	http://en.wikipedia.org/wiki/David_Foster
David Foster Wallace	http://en.wikipedia.org/wiki/David_Foster_Wallace
David Friedrich Strauss	http://en.wikipedia.org/wiki/David_Friedrich_Strauss
David Frost	http://en.wikipedia.org/wiki/David_Frost
David Frum	http://en.wikipedia.org/wiki/David_Frum
David Fuhrer	http://en.wikipedia.org/wiki/David_Fuhrer
David Gallagher	http://en.wikipedia.org/wiki/David_Gallagher
David Garnett	http://en.wikipedia.org/wiki/David_Garnett
David Garrick	http://en.wikipedia.org/wiki/David_Garrick
David Gauke	http://en.wikipedia.org/wiki/David_Gauke
David Geffen	http://en.wikipedia.org/wiki/David_Geffen
David Gergen	http://en.wikipedia.org/wiki/David_Gergen
David Gest	http://en.wikipedia.org/wiki/David_Gest
David Gilmour	http://en.wikipedia.org/wiki/David_Gilmour
David Goodnow	http://en.wikipedia.org/wiki/David_Goodnow
David Graf	http://en.wikipedia.org/wiki/David_Graf
David Graham Phillips	http://en.wikipedia.org/wiki/David_Graham_Phillips
David Greenglass	http://en.wikipedia.org/wiki/David_Greenglass
David Gregory	http://en.wikipedia.org/wiki/David_Gregory_(journalist)
David Grossman	http://en.wikipedia.org/wiki/David_Grossman
David Halberstam	http://en.wikipedia.org/wiki/David_Halberstam
David Hamilton	http://en.wikipedia.org/wiki/David_Hamilton_(politician)
David Hanson	http://en.wikipedia.org/wiki/David_Hanson_(politician)
David Harris	http://en.wikipedia.org/wiki/David_Harris
David Hartley	http://en.wikipedia.org/wiki/David_Hartley_(philosopher)
David Hartman	http://en.wikipedia.org/wiki/David_Hartman_(TV_personality)
David Hasselhoff	http://en.wikipedia.org/wiki/David_Hasselhoff
David Heath	http://en.wikipedia.org/wiki/David_Heath
David Hedison	http://en.wikipedia.org/wiki/David_Hedison
David Helfgott	http://en.wikipedia.org/wiki/David_Helfgott
David Hemmings	http://en.wikipedia.org/wiki/David_Hemmings
David Heyes	http://en.wikipedia.org/wiki/David_Heyes
David Hicks	http://en.wikipedia.org/wiki/David_Hicks
David Hilbert	http://en.wikipedia.org/wiki/David_Hilbert
David Hobson	http://en.wikipedia.org/wiki/Dave_Hobson
David Hockney	http://en.wikipedia.org/wiki/David_Hockney
David Hodo	http://en.wikipedia.org/wiki/David_Hodo
David Hookes	http://en.wikipedia.org/wiki/David_Hookes
David Horowitz	http://en.wikipedia.org/wiki/David_Horowitz
David Huddleston	http://en.wikipedia.org/wiki/David_Huddleston
David Hughes	http://en.wikipedia.org/wiki/David_Hughes_%28musician%29
David Hume	http://en.wikipedia.org/wiki/David_Hume
David Hyde Pierce	http://en.wikipedia.org/wiki/David_Hyde_Pierce
David I	http://en.wikipedia.org/wiki/David_I_of_Scotland
David Icke	http://en.wikipedia.org/wiki/David_Icke
David Ignatow	http://en.wikipedia.org/wiki/David_Ignatow
David II	http://en.wikipedia.org/wiki/David_II
David Irving	http://en.wikipedia.org/wiki/David_Irving
David J. O'Reilly	http://en.wikipedia.org/wiki/David_J._O%27Reilly
David J. Stern	http://en.wikipedia.org/wiki/David_J._Stern
David James Elliott	http://en.wikipedia.org/wiki/David_James_Elliott
David Janssen	http://en.wikipedia.org/wiki/David_Janssen
David Jason	http://en.wikipedia.org/wiki/David_Jason
David Johansen	http://en.wikipedia.org/wiki/David_Johansen
David Jones	http://en.wikipedia.org/wiki/David_Jones_(Welsh_politician)
David Justice	http://en.wikipedia.org/wiki/David_Justice
David K. E. Bruce	http://en.wikipedia.org/wiki/David_K._E._Bruce
David Kay	http://en.wikipedia.org/wiki/David_Kay
David Keene	http://en.wikipedia.org/wiki/David_Keene
David Keith	http://en.wikipedia.org/wiki/David_Keith
David Knopfler	http://en.wikipedia.org/wiki/David_Knopfler
David Koresh	http://en.wikipedia.org/wiki/David_Koresh
David Krumholtz	http://en.wikipedia.org/wiki/David_Krumholtz
David L. Boren	http://en.wikipedia.org/wiki/David_L._Boren
David L. Boren	http://en.wikipedia.org/wiki/David_L._Boren
David L. Clarke	http://en.wikipedia.org/wiki/David_L._Clarke
David L. Lander	http://en.wikipedia.org/wiki/David_L._Lander
David L. Wolper	http://en.wikipedia.org/wiki/David_L._Wolper
David Lammy	http://en.wikipedia.org/wiki/David_Lammy
David Lascher	http://en.wikipedia.org/wiki/David_Lascher
David Laws	http://en.wikipedia.org/wiki/David_Laws
David Lean	http://en.wikipedia.org/wiki/David_Lean
David Leavitt	http://en.wikipedia.org/wiki/David_Leavitt
David Lee Roth	http://en.wikipedia.org/wiki/David_Lee_Roth
David Leisure	http://en.wikipedia.org/wiki/David_Leisure
David Letterman	http://en.wikipedia.org/wiki/David_Letterman
David Lidington	http://en.wikipedia.org/wiki/David_Lidington
David Livingstone	http://en.wikipedia.org/wiki/David_Livingstone
David Lloyd George	http://en.wikipedia.org/wiki/David_Lloyd_George
David Lodge	http://en.wikipedia.org/wiki/David_Lodge_(author)
David Lovering	http://en.wikipedia.org/wiki/David_Lovering
David Lowery	http://en.wikipedia.org/wiki/David_Lowery
David Lynch	http://en.wikipedia.org/wiki/David_Lynch
David M. Halperin	http://en.wikipedia.org/wiki/David_M._Halperin
David M. Lee	http://en.wikipedia.org/wiki/David_M._Lee
David M. Navarro	http://en.wikipedia.org/wiki/Dave_Navarro
David M. Rubenstein	http://en.wikipedia.org/wiki/David_M._Rubenstein
David M. Thomas	http://en.wikipedia.org/wiki/David_M._Thomas
David Mamet	http://en.wikipedia.org/wiki/David_Mamet
David Martin	http://en.wikipedia.org/wiki/David_O'Brien_Martin
David Maysles	http://en.wikipedia.org/wiki/David_Maysles
David McCallum	http://en.wikipedia.org/wiki/David_McCallum
David McCullough	http://en.wikipedia.org/wiki/David_McCullough
David McIntosh	http://en.wikipedia.org/wiki/David_M._McIntosh
David Miliband	http://en.wikipedia.org/wiki/David_Miliband
David Minge	http://en.wikipedia.org/wiki/David_Minge
David Miscavige	http://en.wikipedia.org/wiki/David_Miscavige
David Morris	http://en.wikipedia.org/wiki/David_Morris_(English_politician)
David Morse	http://en.wikipedia.org/wiki/David_Morse_(actor)
David Mowat	http://en.wikipedia.org/wiki/David_Mowat
David Mundell	http://en.wikipedia.org/wiki/David_Mundell
David Narcizo	http://en.wikipedia.org/wiki/David_Narcizo
David Naughton	http://en.wikipedia.org/wiki/David_Naughton_(actor)
David Neeleman	http://en.wikipedia.org/wiki/David_Neeleman
David Nelson	http://en.wikipedia.org/wiki/David_Nelson_(actor)
David Niven	http://en.wikipedia.org/wiki/David_Niven
David Nuttall	http://en.wikipedia.org/wiki/David_Nuttall
David O. Selznick	http://en.wikipedia.org/wiki/David_O._Selznick
David Obey	http://en.wikipedia.org/wiki/David_Obey
David Oddsson	http://en.wikipedia.org/wiki/David_Oddsson
David Ogden Stiers	http://en.wikipedia.org/wiki/David_Ogden_Stiers
David Ortiz	http://en.wikipedia.org/wiki/David_Ortiz
David P. Buckson	http://en.wikipedia.org/wiki/David_P._Buckson
David Pack	http://en.wikipedia.org/wiki/David_Pack
David Packard	http://en.wikipedia.org/wiki/David_Packard
David Palmer	http://en.wikipedia.org/wiki/Dee_Palmer
David Petraeus	http://en.wikipedia.org/wiki/David_Petraeus
David Phelps	http://en.wikipedia.org/wiki/David_Phelps
David Pinski	http://en.wikipedia.org/wiki/David_Pinski
David Pratt	http://en.wikipedia.org/wiki/David_Pratt_(politician)
David Price	http://en.wikipedia.org/wiki/David_Price_(American_politician)
David Proval	http://en.wikipedia.org/wiki/David_Proval
David Prowse	http://en.wikipedia.org/wiki/David_Prowse
David Pryor	http://en.wikipedia.org/wiki/David_Pryor
David Pryor	http://en.wikipedia.org/wiki/David_Pryor
David R. Goode	http://en.wikipedia.org/wiki/David_R._Goode
David R. Obey	http://en.wikipedia.org/wiki/David_R._Obey
David Rabe	http://en.wikipedia.org/wiki/David_Rabe
David Rakoff	http://en.wikipedia.org/wiki/David_Rakoff
David Rees	http://en.wikipedia.org/wiki/David_Rees_(cartoonist)
David Reimer	http://en.wikipedia.org/wiki/David_Reimer
David Remnick	http://en.wikipedia.org/wiki/David_Remnick
David Ricardo	http://en.wikipedia.org/wiki/David_Ricardo
David Rice Atchison	http://en.wikipedia.org/wiki/David_Rice_Atchison
David Robinson	http://en.wikipedia.org/wiki/David_Robinson_(basketball)
David Rockefeller	http://en.wikipedia.org/wiki/David_Rockefeller
David Ruffin	http://en.wikipedia.org/wiki/David_Ruffin
David Ruffley	http://en.wikipedia.org/wiki/David_Ruffley
David Rutley	http://en.wikipedia.org/wiki/David_Rutley
David S. Monson	http://en.wikipedia.org/wiki/David_S._Monson
David Safavian	http://en.wikipedia.org/wiki/David_Safavian
David Sanborn	http://en.wikipedia.org/wiki/David_Sanborn
David Sarnoff	http://en.wikipedia.org/wiki/David_Sarnoff
David Satcher	http://en.wikipedia.org/wiki/David_Satcher
David Schwimmer	http://en.wikipedia.org/wiki/David_Schwimmer
David Scott	http://en.wikipedia.org/wiki/David_Scott_(Georgia)
David Sedaris	http://en.wikipedia.org/wiki/David_Sedaris
David Selby	http://en.wikipedia.org/wiki/David_Selby
David Simon	http://en.wikipedia.org/wiki/David_Simon
David Simon	http://en.wikipedia.org/wiki/David_Simon
David Simpson	http://en.wikipedia.org/wiki/David_Simpson_(UK_politician)
David Skaggs	http://en.wikipedia.org/wiki/David_Skaggs
David Soul	http://en.wikipedia.org/wiki/David_Soul
David Souter	http://en.wikipedia.org/wiki/David_Souter
David Spade	http://en.wikipedia.org/wiki/David_Spade
David Steinberg	http://en.wikipedia.org/wiki/David_Steinberg
David Stockman	http://en.wikipedia.org/wiki/David_Stockman
David Storey	http://en.wikipedia.org/wiki/David_Storey
David Strathairn	http://en.wikipedia.org/wiki/David_Strathairn
David Strickland	http://en.wikipedia.org/wiki/David_Strickland
David Suchet	http://en.wikipedia.org/wiki/David_Suchet
David Sutcliffe	http://en.wikipedia.org/wiki/David_Sutcliffe
David Suzuki	http://en.wikipedia.org/wiki/David_Suzuki
David Sylvian	http://en.wikipedia.org/wiki/David_Sylvian
David T. Kearns	http://en.wikipedia.org/wiki/David_T._Kearns
David Talbot	http://en.wikipedia.org/wiki/David_Talbot
David Teniers the Elder	http://en.wikipedia.org/wiki/David_Teniers_the_Elder
David Teniers the Younger	http://en.wikipedia.org/wiki/David_Teniers_the_Younger
David Tennant	http://en.wikipedia.org/wiki/David_Tennant
David Thewlis	http://en.wikipedia.org/wiki/David_Thewlis
David Thomas	http://en.wikipedia.org/wiki/David_Thomas_(musician)
David Thompson	http://en.wikipedia.org/wiki/David_Thompson_(Barbadian_politician)
David Tibet	http://en.wikipedia.org/wiki/David_Tibet
David Tomlinson	http://en.wikipedia.org/wiki/David_Tomlinson
David Tredinnick	http://en.wikipedia.org/wiki/David_Tredinnick_(politician)
David Trimble	http://en.wikipedia.org/wiki/David_Trimble
David Trimble	http://en.wikipedia.org/wiki/David_Trimble
David Tudor	http://en.wikipedia.org/wiki/David_Tudor
David Urquhart	http://en.wikipedia.org/wiki/David_Urquhart
David Vetter	http://en.wikipedia.org/wiki/David_Vetter
David Vitter	http://en.wikipedia.org/wiki/David_Vitter
David W. Dorman	http://en.wikipedia.org/wiki/David_W._Dorman
David Wain	http://en.wikipedia.org/wiki/David_Wain
David Walliams	http://en.wikipedia.org/wiki/David_Walliams
David Ward	http://en.wikipedia.org/wiki/David_Ward_(politician)
David Warner	http://en.wikipedia.org/wiki/David_Warner_(actor)
David Wells	http://en.wikipedia.org/wiki/David_Wells
David Wenham	http://en.wikipedia.org/wiki/David_Wenham
David White	http://en.wikipedia.org/wiki/David_White_(actor)
David Willetts	http://en.wikipedia.org/wiki/David_Willetts
David Winnick	http://en.wikipedia.org/wiki/David_Winnick
David Wise	http://en.wikipedia.org/wiki/David_Wise_%28writer%29
David Wm Sims	http://en.wikipedia.org/wiki/David_Wm._Sims
David Wright	http://en.wikipedia.org/wiki/David_Wright_(politician)
David Wu	http://en.wikipedia.org/wiki/David_Wu
David X. Cohen	http://en.wikipedia.org/wiki/David_X._Cohen
David Yow	http://en.wikipedia.org/wiki/David_Yow
Davy Crockett	http://en.wikipedia.org/wiki/Davy_Crockett
Davy Jones	http://en.wikipedia.org/wiki/David_Jones_(jazz_musician)
Dawn Fraser	http://en.wikipedia.org/wiki/Dawn_Fraser
Dawn French	http://en.wikipedia.org/wiki/Dawn_French
Dawn McCarthy	http://en.wikipedia.org/wiki/Dawn_McCarthy
Dawn Penn	http://en.wikipedia.org/wiki/Dawn_Penn
Dawn Powell	http://en.wikipedia.org/wiki/Dawn_Powell
Dawn Primarolo	http://en.wikipedia.org/wiki/Dawn_Primarolo
Dawn Wells	http://en.wikipedia.org/wiki/Dawn_Wells
Dayo Ade	http://en.wikipedia.org/wiki/Dayo_Ade
Dayton Leroy Rogers	http://en.wikipedia.org/wiki/Dayton_Leroy_Rogers
Dayyan Eng	http://en.wikipedia.org/wiki/Dayyan_Eng
De Witt Clinton	http://en.wikipedia.org/wiki/De_Witt_Clinton
Deal Hudson	http://en.wikipedia.org/wiki/Deal_Hudson
Dean A. Gallo	http://en.wikipedia.org/wiki/Dean_A._Gallo
Dean Acheson	http://en.wikipedia.org/wiki/Dean_Acheson
Dean Barrow	http://en.wikipedia.org/wiki/Dean_Barrow
Dean Cain	http://en.wikipedia.org/wiki/Dean_Cain
Dean Cameron	http://en.wikipedia.org/wiki/Dean_Cameron
Dean Haglund	http://en.wikipedia.org/wiki/Dean_Haglund
Dean Heller	http://en.wikipedia.org/wiki/Dean_Heller
Dean Jagger	http://en.wikipedia.org/wiki/Dean_Jagger
Dean Jones	http://en.wikipedia.org/wiki/Dean_Jones_(actor)
Dean Jones	http://en.wikipedia.org/wiki/Dean_Jones_(cricketer)
Dean Kamen	http://en.wikipedia.org/wiki/Dean_Kamen
Dean Martin	http://en.wikipedia.org/wiki/Dean_Martin
Dean R. Koontz	http://en.wikipedia.org/wiki/Dean_R._Koontz
Dean Rusk	http://en.wikipedia.org/wiki/Dean_Rusk
Dean Stockwell	http://en.wikipedia.org/wiki/Dean_Stockwell
Dean Torrence	http://en.wikipedia.org/wiki/Dean_Torrence
Dean Ween	http://en.wikipedia.org/wiki/Dean_Ween
Dean Winters	http://en.wikipedia.org/wiki/Dean_Winters
Deanna Durbin	http://en.wikipedia.org/wiki/Deanna_Durbin
Dean-Paul Martin	http://en.wikipedia.org/wiki/Dean_Paul_Martin
Debbi Fields	http://en.wikipedia.org/wiki/Debbi_Fields
Debbi Peterson	http://en.wikipedia.org/wiki/Debbi_Peterson
Debbie Allen	http://en.wikipedia.org/wiki/Debbie_Allen
Debbie Gibson	http://en.wikipedia.org/wiki/Debbie_Gibson
Debbie Halvorson	http://en.wikipedia.org/wiki/Debbie_Halvorson
Debbie Harry	http://en.wikipedia.org/wiki/Debbie_Harry
Debbie Reynolds	http://en.wikipedia.org/wiki/Debbie_Reynolds
Debbie Rowe	http://en.wikipedia.org/wiki/Debbie_Rowe
Debbie Stabenow	http://en.wikipedia.org/wiki/Debbie_Stabenow
Debbie Stoller	http://en.wikipedia.org/wiki/Debbie_Stoller
Debbie Wasserman Schultz	http://en.wikipedia.org/wiki/Debbie_Wasserman_Schultz
Debby Boone	http://en.wikipedia.org/wiki/Debby_Boone
Debi Mazar	http://en.wikipedia.org/wiki/Debi_Mazar
Deborah Bull	http://en.wikipedia.org/wiki/Deborah_Bull
Deborah Harry	http://en.wikipedia.org/wiki/Deborah_Harry
Deborah Jin	http://en.wikipedia.org/wiki/Deborah_Jin
Deborah Kerr	http://en.wikipedia.org/wiki/Deborah_Kerr
Deborah Norville	http://en.wikipedia.org/wiki/Deborah_Norville
Deborah Pryce	http://en.wikipedia.org/wiki/Deborah_Pryce
Deborah Raffin	http://en.wikipedia.org/wiki/Deborah_Raffin
Deborah Tannen	http://en.wikipedia.org/wiki/Deborah_Tannen
Deborah Walley	http://en.wikipedia.org/wiki/Deborah_Walley
Debra Byrd	http://en.wikipedia.org/wiki/Debra_Byrd
Debra Jo Rupp	http://en.wikipedia.org/wiki/Debra_Jo_Rupp
Debra Messing	http://en.wikipedia.org/wiki/Debra_Messing
Debra Paget	http://en.wikipedia.org/wiki/Debra_Paget
Debra Wasserman	http://en.wikipedia.org/wiki/Debbie_Wasserman_Schultz
Debra Wilson	http://en.wikipedia.org/wiki/Debra_Wilson
Debra Winger	http://en.wikipedia.org/wiki/Debra_Winger
Debralee Scott	http://en.wikipedia.org/wiki/Debralee_Scott
Declan McCullagh	http://en.wikipedia.org/wiki/Declan_McCullagh
Dede Allen	http://en.wikipedia.org/wiki/Dede_Allen
Dedee Pfeiffer	http://en.wikipedia.org/wiki/Dedee_Pfeiffer
Dee Dee Myers	http://en.wikipedia.org/wiki/Dee_Dee_Myers
Dee Dee Ramone	http://en.wikipedia.org/wiki/Dee_Dee_Ramone
Dee Dee Warwick	http://en.wikipedia.org/wiki/Dee_Dee_Warwick
Dee Snider	http://en.wikipedia.org/wiki/Dee_Snider
Dee Wallace-Stone	http://en.wikipedia.org/wiki/Dee_Wallace-Stone
Deep Roy	http://en.wikipedia.org/wiki/Deep_Roy
Deepak Chopra	http://en.wikipedia.org/wiki/Deepak_Chopra
DeForest Kelley	http://en.wikipedia.org/wiki/DeForest_Kelley
DeForest Soaries	http://en.wikipedia.org/wiki/DeForest_Soaries
Deidre Hall	http://en.wikipedia.org/wiki/Deidre_Hall
Deion Sanders	http://en.wikipedia.org/wiki/Deion_Sanders
Del Shannon	http://en.wikipedia.org/wiki/Del_Shannon
Del Tha Funkee Homosapien	http://en.wikipedia.org/wiki/Del_Tha_Funkee_Homosapien
Delaney Williams	http://en.wikipedia.org/wiki/Delaney_Williams
Delbert L. Latta	http://en.wikipedia.org/wiki/Delbert_L._Latta
Delbert Mann	http://en.wikipedia.org/wiki/Delbert_Mann
Delia Bacon	http://en.wikipedia.org/wiki/Delia_Bacon
Delia Derbyshire	http://en.wikipedia.org/wiki/Delia_Derbyshire
Della Reese	http://en.wikipedia.org/wiki/Della_Reese
Delmer Daves	http://en.wikipedia.org/wiki/Delmer_Daves
Delmore Schwartz	http://en.wikipedia.org/wiki/Delmore_Schwartz
Delroy Lindo	http://en.wikipedia.org/wiki/Delroy_Lindo
Delta Burke	http://en.wikipedia.org/wiki/Delta_Burke
Delta Goodrem	http://en.wikipedia.org/wiki/Delta_Goodrem
Demi Moore	http://en.wikipedia.org/wiki/Demi_Moore
Demond Wilson	http://en.wikipedia.org/wiki/Demond_Wilson
Denardo Coleman	http://en.wikipedia.org/wiki/Denardo_Coleman
Deng Xiaoping	http://en.wikipedia.org/wiki/Deng_Xiaoping
Denholm Elliott	http://en.wikipedia.org/wiki/Denholm_Elliott
Deniece Williams	http://en.wikipedia.org/wiki/Deniece_Williams
Denis Diderot	http://en.wikipedia.org/wiki/Denis_Diderot
Denis Johnson	http://en.wikipedia.org/wiki/Denis_Johnson
Denis Law	http://en.wikipedia.org/wiki/Denis_Law
Denis Leary	http://en.wikipedia.org/wiki/Denis_Leary
Denis Mackail	http://en.wikipedia.org/wiki/Denis_Mackail
Denis MacShane	http://en.wikipedia.org/wiki/Denis_MacShane
Denis Papin	http://en.wikipedia.org/wiki/Denis_Papin
Denis Sassou-Nguesso	http://en.wikipedia.org/wiki/Denis_Sassou-Nguesso
Denise Black	http://en.wikipedia.org/wiki/Denise_Black
Denise Crosby	http://en.wikipedia.org/wiki/Denise_Crosby
Denise Levertov	http://en.wikipedia.org/wiki/Denise_Levertov
Denise Majette	http://en.wikipedia.org/wiki/Denise_Majette
Denise Rich	http://en.wikipedia.org/wiki/Denise_Rich
Denise Richards	http://en.wikipedia.org/wiki/Denise_Richards
Denise van Outen	http://en.wikipedia.org/wiki/Denise_van_Outen
Denise Welch	http://en.wikipedia.org/wiki/Denise_Welch
Dennis Bergkamp	http://en.wikipedia.org/wiki/Dennis_Bergkamp
Dennis Brutus	http://en.wikipedia.org/wiki/Dennis_Brutus
Dennis Cardoza	http://en.wikipedia.org/wiki/Dennis_Cardoza
Dennis Christopher	http://en.wikipedia.org/wiki/Dennis_Christopher
Dennis Crosby	http://en.wikipedia.org/wiki/Dennis_Crosby
Dennis Day	http://en.wikipedia.org/wiki/Dennis_Day
Dennis DeConcini	http://en.wikipedia.org/wiki/Dennis_DeConcini
Dennis DeConcini	http://en.wikipedia.org/wiki/Dennis_DeConcini
Dennis Dugan	http://en.wikipedia.org/wiki/Dennis_Dugan
Dennis E. Eckart	http://en.wikipedia.org/wiki/Dennis_E._Eckart
Dennis Eckersley	http://en.wikipedia.org/wiki/Dennis_Eckersley
Dennis Erectus	http://en.wikipedia.org/wiki/Dennis_Erectus
Dennis Farina	http://en.wikipedia.org/wiki/Dennis_Farina
Dennis Franz	http://en.wikipedia.org/wiki/Dennis_Franz
Dennis Gabor	http://en.wikipedia.org/wiki/Dennis_Gabor
Dennis Hastert	http://en.wikipedia.org/wiki/Dennis_Hastert
Dennis Haysbert	http://en.wikipedia.org/wiki/Dennis_Haysbert
Dennis Hopper	http://en.wikipedia.org/wiki/Dennis_Hopper
Dennis Kozlowski	http://en.wikipedia.org/wiki/Dennis_Kozlowski
Dennis Kucinich	http://en.wikipedia.org/wiki/Dennis_Kucinich
Dennis Kucinich	http://en.wikipedia.org/wiki/Dennis_Kucinich
Dennis M. Hertel	http://en.wikipedia.org/wiki/Dennis_M._Hertel
Dennis Miller	http://en.wikipedia.org/wiki/Dennis_Miller
Dennis Moore	http://en.wikipedia.org/wiki/Dennis_Moore
Dennis Morgan	http://en.wikipedia.org/wiki/Dennis_Morgan
Dennis Muren	http://en.wikipedia.org/wiki/Dennis_Muren
Dennis Prager	http://en.wikipedia.org/wiki/Dennis_Prager
Dennis Quaid	http://en.wikipedia.org/wiki/Dennis_Quaid
Dennis Rader	http://en.wikipedia.org/wiki/Dennis_Rader
Dennis Rehberg	http://en.wikipedia.org/wiki/Dennis_Rehberg
Dennis Ritchie	http://en.wikipedia.org/wiki/Dennis_Ritchie
Dennis Rodman	http://en.wikipedia.org/wiki/Dennis_Rodman
Dennis Skinner	http://en.wikipedia.org/wiki/Dennis_Skinner
Dennis Weaver	http://en.wikipedia.org/wiki/Dennis_Weaver
Dennis Weaver	http://en.wikipedia.org/wiki/Dennis_Weaver
Dennis Wilson	http://en.wikipedia.org/wiki/Dennis_Wilson
Denny Laine	http://en.wikipedia.org/wiki/Denny_Laine
Denny McLain	http://en.wikipedia.org/wiki/Denny_McLain
Denny Seiwell	http://en.wikipedia.org/wiki/Denny_Seiwell
Denny Smith	http://en.wikipedia.org/wiki/Denny_Smith
Denver Pyle	http://en.wikipedia.org/wiki/Denver_Pyle
Denys Lasdun	http://en.wikipedia.org/wiki/Denys_Lasdun
Denzel Washington	http://en.wikipedia.org/wiki/Denzel_Washington
Denzil Douglas	http://en.wikipedia.org/wiki/Denzil_Douglas
Deodoro da Fonseca	http://en.wikipedia.org/wiki/Deodoro_da_Fonseca
Derek Bailey	http://en.wikipedia.org/wiki/Derek_Bailey
Derek Barton	http://en.wikipedia.org/wiki/Derek_Barton
Derek Bok	http://en.wikipedia.org/wiki/Derek_Bok
Derek Jacobi	http://en.wikipedia.org/wiki/Derek_Jacobi
Derek Jarman	http://en.wikipedia.org/wiki/Derek_Jarman
Derek Jeter	http://en.wikipedia.org/wiki/Derek_Jeter
Derek Mahon	http://en.wikipedia.org/wiki/Derek_Mahon
Derek Sikua	http://en.wikipedia.org/wiki/Derek_Sikua
Derek Twigg	http://en.wikipedia.org/wiki/Derek_Twigg
Derek Walcott	http://en.wikipedia.org/wiki/Derek_Walcott
Dermot Mulroney	http://en.wikipedia.org/wiki/Dermot_Mulroney
Derya Alabora	http://en.wikipedia.org/wiki/Derya_Alabora
Deryck Whibley	http://en.wikipedia.org/wiki/Deryck_Whibley
Des McAnuff	http://en.wikipedia.org/wiki/Des_McAnuff
DeShaun Holton	http://en.wikipedia.org/wiki/DeShaun_Holton
Desi Arnaz	http://en.wikipedia.org/wiki/Desi_Arnaz
Desi Arnaz, Jr.	http://en.wikipedia.org/wiki/Desi_Arnaz%2C_Jr.
Desiderio da Settignano	http://en.wikipedia.org/wiki/Desiderio_da_Settignano
Desmond Dekker	http://en.wikipedia.org/wiki/Desmond_Dekker
Desmond Harrington	http://en.wikipedia.org/wiki/Desmond_Harrington
Desmond Howard	http://en.wikipedia.org/wiki/Desmond_Howard
Desmond Llewelyn	http://en.wikipedia.org/wiki/Desmond_Llewelyn
Desmond Swayne	http://en.wikipedia.org/wiki/Desmond_Swayne
Desmond Tutu	http://en.wikipedia.org/wiki/Desmond_Tutu
Devendra Banhart	http://en.wikipedia.org/wiki/Devendra_Banhart
Devin Nunes	http://en.wikipedia.org/wiki/Devin_Nunes
Devon Aoki	http://en.wikipedia.org/wiki/Devon_Aoki
Devon Sawa	http://en.wikipedia.org/wiki/Devon_Sawa
Devon Scott	http://en.wikipedia.org/wiki/Devon_Scott
Dewey Bunnell	http://en.wikipedia.org/wiki/Dewey_Bunnell
DeWitt Wallace	http://en.wikipedia.org/wiki/DeWitt_Wallace
Dexter Fletcher	http://en.wikipedia.org/wiki/Dexter_Fletcher
Dexter Holland	http://en.wikipedia.org/wiki/Dexter_Holland
Diahann Carroll	http://en.wikipedia.org/wiki/Diahann_Carroll
Dian Fossey	http://en.wikipedia.org/wiki/Dian_Fossey
Diana DeGette	http://en.wikipedia.org/wiki/Diana_DeGette
Diana Dors	http://en.wikipedia.org/wiki/Diana_Dors
Diana Hyland	http://en.wikipedia.org/wiki/Diana_Hyland
Diana Krall	http://en.wikipedia.org/wiki/Diana_Krall
Diana Lynn	http://en.wikipedia.org/wiki/Diana_Lynn
Diana Muldaur	http://en.wikipedia.org/wiki/Diana_Muldaur
Diana R. Johnson	http://en.wikipedia.org/wiki/Diana_Johnson
Diana Rigg	http://en.wikipedia.org/wiki/Diana_Rigg
Diana Ross	http://en.wikipedia.org/wiki/Diana_Ross
Diana Trilling	http://en.wikipedia.org/wiki/Diana_Trilling
Diane Abbott	http://en.wikipedia.org/wiki/Diane_Abbott
Diane Ackerman	http://en.wikipedia.org/wiki/Diane_Ackerman
Diane Arbus	http://en.wikipedia.org/wiki/Diane_Arbus
Diane de France	http://en.wikipedia.org/wiki/Diane_de_France
Diane de Poitiers	http://en.wikipedia.org/wiki/Diane_de_Poitiers
Diane Johnson	http://en.wikipedia.org/wiki/Diane_Johnson
Diane Keaton	http://en.wikipedia.org/wiki/Diane_Keaton
Diane Kruger	http://en.wikipedia.org/wiki/Diane_Kruger
Diane Ladd	http://en.wikipedia.org/wiki/Diane_Ladd
Diane Lane	http://en.wikipedia.org/wiki/Diane_Lane
Diane McBain	http://en.wikipedia.org/wiki/Diane_McBain
Diane Neal	http://en.wikipedia.org/wiki/Diane_Neal
Diane Ravitch	http://en.wikipedia.org/wiki/Diane_Ravitch
Diane Sawyer	http://en.wikipedia.org/wiki/Diane_Sawyer
Diane Schuur	http://en.wikipedia.org/wiki/Diane_Schuur
Diane von Furstenberg	http://en.wikipedia.org/wiki/Diane_von_Furstenberg
Diane Wakoski	http://en.wikipedia.org/wiki/Diane_Wakoski
Diane Watson	http://en.wikipedia.org/wiki/Diane_Watson
Dianne Feinstein	http://en.wikipedia.org/wiki/Dianne_Feinstein
Dianne Wiest	http://en.wikipedia.org/wiki/Dianne_Wiest
Dick Armey	http://en.wikipedia.org/wiki/Dick_Armey
Dick Butkus	http://en.wikipedia.org/wiki/Dick_Butkus
Dick Button	http://en.wikipedia.org/wiki/Dick_Button
Dick Cavett	http://en.wikipedia.org/wiki/Dick_Cavett
Dick Cheney	http://en.wikipedia.org/wiki/Dick_Cheney
Dick Cheney	http://en.wikipedia.org/wiki/Dick_Cheney
Dick Clark	http://en.wikipedia.org/wiki/Dick_Clark
Dick Dale	http://en.wikipedia.org/wiki/Dick_Dale
Dick Durbin	http://en.wikipedia.org/wiki/Dick_Durbin
Dick Ebersol	http://en.wikipedia.org/wiki/Dick_Ebersol
Dick Fosbury	http://en.wikipedia.org/wiki/Dick_Fosbury
Dick Francis	http://en.wikipedia.org/wiki/Dick_Francis
Dick Gautier	http://en.wikipedia.org/wiki/Dick_Gautier
Dick Gephardt	http://en.wikipedia.org/wiki/Dick_Gephardt
Dick Gregory	http://en.wikipedia.org/wiki/Dick_Gregory
Dick Haymes	http://en.wikipedia.org/wiki/Dick_Haymes
Dick Hyman	http://en.wikipedia.org/wiki/Dick_Hyman
Dick Lugar	http://en.wikipedia.org/wiki/Dick_Lugar
Dick Martin	http://en.wikipedia.org/wiki/Dick_Martin_(comedian)
Dick Morris	http://en.wikipedia.org/wiki/Dick_Morris
Dick Mountjoy	http://en.wikipedia.org/wiki/Dick_Mountjoy
Dick Powell	http://en.wikipedia.org/wiki/Dick_Powell
Dick Riordan	http://en.wikipedia.org/wiki/Dick_Riordan
Dick Sargent	http://en.wikipedia.org/wiki/Dick_Sargent
Dick Schaap	http://en.wikipedia.org/wiki/Dick_Schaap
Dick Schulze	http://en.wikipedia.org/wiki/Dick_Schulze
Dick Shawn	http://en.wikipedia.org/wiki/Dick_Shawn
Dick Smothers	http://en.wikipedia.org/wiki/Dick_Smothers
Dick Thornburgh	http://en.wikipedia.org/wiki/Dick_Thornburgh
Dick Trickle	http://en.wikipedia.org/wiki/Dick_Trickle
Dick Turpin	http://en.wikipedia.org/wiki/Dick_Turpin
Dick Van Dyke	http://en.wikipedia.org/wiki/Dick_Van_Dyke
Dick Van Patten	http://en.wikipedia.org/wiki/Dick_Van_Patten
Dick Vitale	http://en.wikipedia.org/wiki/Dick_Vitale
Dick Weber	http://en.wikipedia.org/wiki/Dick_Weber
Dick Whittington	http://en.wikipedia.org/wiki/Dick_Whittington
Dick Wolf	http://en.wikipedia.org/wiki/Dick_Wolf
Dick York	http://en.wikipedia.org/wiki/Dick_York
Dickie Bird	http://en.wikipedia.org/wiki/Dickie_Bird
Dickie Jones	http://en.wikipedia.org/wiki/Dickie_Jones
Dickie Moore	http://en.wikipedia.org/wiki/Dickie_Moore_(actor)
Didius Julianus	http://en.wikipedia.org/wiki/Didius_Julianus
Diego Abatantuono	http://en.wikipedia.org/wiki/Diego_Abatantuono
Diego Luna	http://en.wikipedia.org/wiki/Diego_Luna
Diego Maradona	http://en.wikipedia.org/wiki/Diego_Maradona
Diego Rivera	http://en.wikipedia.org/wiki/Diego_Rivera
Diego Vel�zquez	http://en.wikipedia.org/wiki/Diego_Vel%C3%A1zquez
Dietrich Buxtehude	http://en.wikipedia.org/wiki/Dietrich_Buxtehude
Dietrich Eckart	http://en.wikipedia.org/wiki/Dietrich_Eckart
Dileita Mohamed Dileita	http://en.wikipedia.org/wiki/Dileita_Mohamed_Dileita
Dillon Anderson	http://en.wikipedia.org/wiki/Dillon_Anderson
Dimebag Darrell	http://en.wikipedia.org/wiki/Dimebag_Darrell
Dimitri from Paris	http://en.wikipedia.org/wiki/Dimitri_from_Paris
Dimitris Christofias	http://en.wikipedia.org/wiki/Dimitris_Christofias
Dina Merrill	http://en.wikipedia.org/wiki/Dina_Merrill
Dina Meyer	http://en.wikipedia.org/wiki/Dina_Meyer
Dina Titus	http://en.wikipedia.org/wiki/Dina_Titus
Dinah Manoff	http://en.wikipedia.org/wiki/Dinah_Manoff
Dinah Sheridan	http://en.wikipedia.org/wiki/Dinah_Sheridan
Dinah Shore	http://en.wikipedia.org/wiki/Dinah_Shore
Dinah Washington	http://en.wikipedia.org/wiki/Dinah_Washington
Dinesh D'Souza	http://en.wikipedia.org/wiki/Dinesh_D%27Souza
Dinmukhammed Akhimov	http://en.wikipedia.org/wiki/Dinmukhammed_Akhimov
Dino De Laurentiis	http://en.wikipedia.org/wiki/Dino_De_Laurentiis
Diogenes La�rtius	http://en.wikipedia.org/wiki/Diogenes_La%C3%Abrtius
Dion Boucicault	http://en.wikipedia.org/wiki/Dion_Boucicault
Dionne Warwick	http://en.wikipedia.org/wiki/Dionne_Warwick
Dionysius Cato	http://en.wikipedia.org/wiki/Dionysius_Cato
Dionysius Exiguus	http://en.wikipedia.org/wiki/Dionysius_Cato
Dionysius Halicarnassus	http://en.wikipedia.org/wiki/Dionysius_Halicarnassus
Dionysius Petavius	http://en.wikipedia.org/wiki/Dionysius_Petavius
Dionysius the Elder	http://en.wikipedia.org/wiki/Dionysius_Thrax
Dionysius the Younger	http://en.wikipedia.org/wiki/Dionysius_Thrax
Dionysius Thrax	http://en.wikipedia.org/wiki/Dionysius_Thrax
Diosdado Macapagal	http://en.wikipedia.org/wiki/Diosdado_Macapagal
Dirk Benedict	http://en.wikipedia.org/wiki/Dirk_Benedict
Dirk Bogarde	http://en.wikipedia.org/wiki/Dirk_Bogarde
Dirk Kempthorne	http://en.wikipedia.org/wiki/Dirk_Kempthorne
Dita Von Teese	http://en.wikipedia.org/wiki/Dita_Von_Teese
Dith Pran	http://en.wikipedia.org/wiki/Dith_Pran
Diva Muffin Zappa	http://en.wikipedia.org/wiki/Diva_Muffin_Zappa
Divine Brown	http://en.wikipedia.org/wiki/Estella_Marie_Thompson
Dixie Carter	http://en.wikipedia.org/wiki/Dixie_Carter
Dixie Dean	http://en.wikipedia.org/wiki/Dixie_Dean
Dixie Lee	http://en.wikipedia.org/wiki/Dixie_Lee
Dixon Denham	http://en.wikipedia.org/wiki/Dixon_Denham
Dizzee Rascal	http://en.wikipedia.org/wiki/Dizzee_Rascal
Dizzy Dean	http://en.wikipedia.org/wiki/Dizzy_Dean
Dizzy Gillespie	http://en.wikipedia.org/wiki/Dizzy_Gillespie
DJ Clue	http://en.wikipedia.org/wiki/DJ_Clue
DJ Danger Mouse	http://en.wikipedia.org/wiki/DJ_Danger_Mouse
DJ Honda	http://en.wikipedia.org/wiki/DJ_Honda
DJ Jazzy Jeff	http://en.wikipedia.org/wiki/DJ_Jazzy_Jeff
DJ Muggs	http://en.wikipedia.org/wiki/DJ_Muggs
DJ Olive	http://en.wikipedia.org/wiki/DJ_Olive
DJ Premier	http://en.wikipedia.org/wiki/DJ_Premier
DJ Qualls	http://en.wikipedia.org/wiki/DJ_Qualls
DJ Quik	http://en.wikipedia.org/wiki/DJ_Quik
DJ Screw	http://en.wikipedia.org/wiki/DJ_Screw
DJ Shadow	http://en.wikipedia.org/wiki/DJ_Shadow
DJ Spooky	http://en.wikipedia.org/wiki/DJ_Spooky
Django Reinhardt	http://en.wikipedia.org/wiki/Django_Reinhardt
Djimon Hounsou	http://en.wikipedia.org/wiki/Djimon_Hounsou
Djuna Barnes	http://en.wikipedia.org/wiki/Djuna_Barnes
Dmitri Mendeleev	http://en.wikipedia.org/wiki/Dmitri_Mendeleev
Dmitri Shostakovich	http://en.wikipedia.org/wiki/Dmitri_Shostakovich
Dmitry Medvedev	http://en.wikipedia.org/wiki/Dmitry_Medvedev
Doc Hastings	http://en.wikipedia.org/wiki/Doc_Hastings
Doc Severinsen	http://en.wikipedia.org/wiki/Doc_Severinsen
Doc Watson	http://en.wikipedia.org/wiki/Doc_Watson
Dodi al-Fayed	http://en.wikipedia.org/wiki/Dodi_al-Fayed
Dog Chapman	http://en.wikipedia.org/wiki/Dog_Chapman
Dolly Parton	http://en.wikipedia.org/wiki/Dolly_Parton
Dolly the sheep	http://en.wikipedia.org/wiki/Dolly_the_sheep
Dolores del Rio	http://en.wikipedia.org/wiki/Dolores_del_Rio
Dolores Hope	http://en.wikipedia.org/wiki/Dolores_Hope
Dolph Lundgren	http://en.wikipedia.org/wiki/Dolph_Lundgren
Dom DeLuise	http://en.wikipedia.org/wiki/Dom_DeLuise
Domenico Cimarosa	http://en.wikipedia.org/wiki/Domenico_Cimarosa
Domenico Ghirlandaio	http://en.wikipedia.org/wiki/Domenico_Ghirlandaio
Domenico Scarlatti	http://en.wikipedia.org/wiki/Domenico_Scarlatti
Dominic Behan	http://en.wikipedia.org/wiki/Dominic_Behan
Dominic Chianese	http://en.wikipedia.org/wiki/Dominic_Chianese
Dominic Grieve	http://en.wikipedia.org/wiki/Dominic_Grieve
Dominic Monaghan	http://en.wikipedia.org/wiki/Dominic_Monaghan
Dominic Purcell	http://en.wikipedia.org/wiki/Dominic_Purcell
Dominic Raab	http://en.wikipedia.org/wiki/Dominic_Raab
Dominic West	http://en.wikipedia.org/wiki/Dominic_West
Dominique A.	http://en.wikipedia.org/wiki/Dominique_A
Dominique de Villepin	http://en.wikipedia.org/wiki/Dominique_de_Villepin
Dominique de Villepin	http://en.wikipedia.org/wiki/Dominique_de_Villepin
Dominique Dunne	http://en.wikipedia.org/wiki/Dominique_Dunne
Dominique Swain	http://en.wikipedia.org/wiki/Dominique_Swain
Dominique Vivant, Baron Denon	http://en.wikipedia.org/wiki/Dominique_Vivant%2C_Baron_Denon
Domino Harvey	http://en.wikipedia.org/wiki/Domino_Harvey
Don Abney	http://en.wikipedia.org/wiki/Don_Abney
Don Adams	http://en.wikipedia.org/wiki/Don_Adams
Don Ameche	http://en.wikipedia.org/wiki/Don_Ameche
Don Amendolia	http://en.wikipedia.org/wiki/Don_Amendolia
Don Bluth	http://en.wikipedia.org/wiki/Don_Bluth
Don Bonker	http://en.wikipedia.org/wiki/Don_Bonker
Don Bradman	http://en.wikipedia.org/wiki/Don_Bradman
Don Callander	http://en.wikipedia.org/wiki/Don_Callander
Don Carcieri	http://en.wikipedia.org/wiki/Don_Carcieri
Don Carlos Buell	http://en.wikipedia.org/wiki/Don_Carlos_Buell
Don Cheadle	http://en.wikipedia.org/wiki/Don_Cheadle
Don Cherry	http://en.wikipedia.org/wiki/Don_Cherry
Don Cornell	http://en.wikipedia.org/wiki/Don_Cornell
Don DeLillo	http://en.wikipedia.org/wiki/Don_DeLillo
Don Dokken	http://en.wikipedia.org/wiki/Don_Dokken
Don Drysdale	http://en.wikipedia.org/wiki/Don_Drysdale
Don Edwards	http://en.wikipedia.org/wiki/Don_Edwards
Don Edwards	http://en.wikipedia.org/wiki/Don_Edwards
Don Everly	http://en.wikipedia.org/wiki/Don_Everly
Don Foster	http://en.wikipedia.org/wiki/Don_Foster_(politician)
Don Fuqua	http://en.wikipedia.org/wiki/Don_Fuqua
Don Gibson	http://en.wikipedia.org/wiki/Don_Gibson
Don Henley	http://en.wikipedia.org/wiki/Don_Henley
Don Herbert	http://en.wikipedia.org/wiki/Don_Herbert
Don Hewitt	http://en.wikipedia.org/wiki/Don_Hewitt
Don Ho	http://en.wikipedia.org/wiki/Don_Ho
Don Imus	http://en.wikipedia.org/wiki/Don_Imus
Don John of Austria	http://en.wikipedia.org/wiki/Don_John_of_Austria
Don John the Younger	http://en.wikipedia.org/wiki/John_of_Austria_the_Younger
Don Johnson	http://en.wikipedia.org/wiki/Don_Johnson
Don King	http://en.wikipedia.org/wiki/Don_King_(boxing_promoter)
Don Kirshner	http://en.wikipedia.org/wiki/Don_Kirshner
Don Knotts	http://en.wikipedia.org/wiki/Don_Knotts
Don LaFontaine	http://en.wikipedia.org/wiki/Don_LaFontaine
Don Larsen	http://en.wikipedia.org/wiki/Don_Larsen
Don Marquis	http://en.wikipedia.org/wiki/Don_Marquis
Don Mattingly	http://en.wikipedia.org/wiki/Don_Mattingly
Don McLean	http://en.wikipedia.org/wiki/Don_McLean
Don Meredith	http://en.wikipedia.org/wiki/Don_Meredith
Don Murphy	http://en.wikipedia.org/wiki/Don_Murphy
Don Nickles	http://en.wikipedia.org/wiki/Don_Nickles
Don Nickles	http://en.wikipedia.org/wiki/Don_Nickles
Don Novello	http://en.wikipedia.org/wiki/Don_Novello
Don Ohlmeyer	http://en.wikipedia.org/wiki/Don_Ohlmeyer
Don Omar	http://en.wikipedia.org/wiki/Don_Omar
Don Pardo	http://en.wikipedia.org/wiki/Don_Pardo
Don Porter	http://en.wikipedia.org/wiki/Don_Porter
Don Preston	http://en.wikipedia.org/wiki/Don_Preston
Don Rickles	http://en.wikipedia.org/wiki/Don_Rickles
Don Riegle	http://en.wikipedia.org/wiki/Don_Riegle
Don Ritter	http://en.wikipedia.org/wiki/Donald_L._Ritter
Don Sherwood	http://en.wikipedia.org/wiki/Don_Sherwood
Don Shula	http://en.wikipedia.org/wiki/Don_Shula
Don Siegel	http://en.wikipedia.org/wiki/Don_Siegel
Don Stark	http://en.wikipedia.org/wiki/Don_Stark
Don Stroud	http://en.wikipedia.org/wiki/Don_Stroud
Don Sundquist	http://en.wikipedia.org/wiki/Don_Sundquist
Don Was	http://en.wikipedia.org/wiki/Don_Was
Don Wildmon	http://en.wikipedia.org/wiki/Don_Wildmon
Don Young	http://en.wikipedia.org/wiki/Don_Young
Don Young	http://en.wikipedia.org/wiki/Don_Young
Don Zimmer	http://en.wikipedia.org/wiki/Don_Zimmer
Donal Logue	http://en.wikipedia.org/wiki/Donal_Logue
Donal Logue	http://en.wikipedia.org/wiki/Donal_Logue
Donald A. Glaser	http://en.wikipedia.org/wiki/Donald_A._Glaser
Donald Barthelme	http://en.wikipedia.org/wiki/Donald_Barthelme
Donald Carcieri	http://en.wikipedia.org/wiki/Donald_Carcieri
Donald Crisp	http://en.wikipedia.org/wiki/Donald_Crisp
Donald Davidson	http://en.wikipedia.org/wiki/Donald_Davidson_(philosopher)
Donald Davidson	http://en.wikipedia.org/wiki/Donald_Davidson_(poet)
Donald E. Graham	http://en.wikipedia.org/wiki/Donald_E._Graham
Donald E. Knuth	http://en.wikipedia.org/wiki/Donald_E._Knuth
Donald Evans	http://en.wikipedia.org/wiki/Donald_Evans
Donald Fagen	http://en.wikipedia.org/wiki/Donald_Fagen
Donald Faison	http://en.wikipedia.org/wiki/Donald_Faison
Donald Gelling	http://en.wikipedia.org/wiki/Donald_Gelling
Donald Grant Mitchell	http://en.wikipedia.org/wiki/Donald_Grant_Mitchell
Donald Hall	http://en.wikipedia.org/wiki/Donald_Hall
Donald Hodel	http://en.wikipedia.org/wiki/Donald_Hodel
Donald J. Carty	http://en.wikipedia.org/wiki/Donald_J._Carty
Donald J. Cram	http://en.wikipedia.org/wiki/Donald_J._Cram
Donald J. Pease	http://en.wikipedia.org/wiki/Donald_J._Pease
Donald James Leslie	http://en.wikipedia.org/wiki/Donald_Leslie
Donald Johanson	http://en.wikipedia.org/wiki/Donald_Johanson
Donald Justice	http://en.wikipedia.org/wiki/Donald_Justice
Donald MacBride	http://en.wikipedia.org/wiki/Donald_MacBride
Donald Manzullo	http://en.wikipedia.org/wiki/Donald_Manzullo
Donald Marron	http://en.wikipedia.org/wiki/Donald_Marron
Donald O'Connor	http://en.wikipedia.org/wiki/Donald_O%27Connor
Donald Ogden Stewart	http://en.wikipedia.org/wiki/Donald_Ogden_Stewart
Donald P. Bellisario	http://en.wikipedia.org/wiki/Donald_P._Bellisario
Donald Payne	http://en.wikipedia.org/wiki/Donald_M._Payne
Donald Petrie	http://en.wikipedia.org/wiki/Donald_Petrie
Donald Pleasence	http://en.wikipedia.org/wiki/Donald_Pleasence
Donald Regan	http://en.wikipedia.org/wiki/Donald_Regan
Donald Rumsfeld	http://en.wikipedia.org/wiki/Donald_Rumsfeld
Donald Segretti	http://en.wikipedia.org/wiki/Donald_Segretti
Donald Sinden	http://en.wikipedia.org/wiki/Donald_Sinden
Donald Sutherland	http://en.wikipedia.org/wiki/Donald_Sutherland
Donald Trump	http://en.wikipedia.org/wiki/Donald_Trump
Donald Tsang	http://en.wikipedia.org/wiki/Donald_Tsang
Donald Tusk	http://en.wikipedia.org/wiki/Donald_Tusk
Donald W. Riegle, Jr.	http://en.wikipedia.org/wiki/Donald_W._Riegle%2C_Jr.
Donatella Versace	http://en.wikipedia.org/wiki/Donatella_Versace
Donato Bramante	http://en.wikipedia.org/wiki/Donato_Bramante
Donna Brazile	http://en.wikipedia.org/wiki/Donna_Brazile
Donna D'Errico	http://en.wikipedia.org/wiki/Donna_D%27Errico
Donna Dixon	http://en.wikipedia.org/wiki/Donna_Dixon
Donna Douglas	http://en.wikipedia.org/wiki/Donna_Douglas
Donna Edwards	http://en.wikipedia.org/wiki/Donna_Edwards
Donna Karan	http://en.wikipedia.org/wiki/Donna_Karan
Donna M. Christian-Christensen	http://en.wikipedia.org/wiki/Donna_M._Christian-Christensen
Donna Mills	http://en.wikipedia.org/wiki/Donna_Mills
Donna Pescow	http://en.wikipedia.org/wiki/Donna_Pescow
Donna Reed	http://en.wikipedia.org/wiki/Donna_Reed
Donna Rice	http://en.wikipedia.org/wiki/Donna_Rice
Donna Shalala	http://en.wikipedia.org/wiki/Donna_Shalala
Donna Summer	http://en.wikipedia.org/wiki/Donna_Summer
Donnie Iris	http://en.wikipedia.org/wiki/Donnie_Iris
Donnie Wahlberg	http://en.wikipedia.org/wiki/Donnie_Wahlberg
Donny Most	http://en.wikipedia.org/wiki/Donny_Most
Donny Osmond	http://en.wikipedia.org/wiki/Donny_Osmond
Donovan McNabb	http://en.wikipedia.org/wiki/Donovan_McNabb
Donovan Scott	http://en.wikipedia.org/wiki/Donovan_Scott
Dontrelle Willis	http://en.wikipedia.org/wiki/Dontrelle_Willis
Doreen Tracey	http://en.wikipedia.org/wiki/Doreen_Tracey
Doris Day	http://en.wikipedia.org/wiki/Doris_Day
Doris Dowling	http://en.wikipedia.org/wiki/Doris_Dowling
Doris Kearns Goodwin	http://en.wikipedia.org/wiki/Doris_Kearns_Goodwin
Doris Kenyon	http://en.wikipedia.org/wiki/Doris_Kenyon
Doris Lessing	http://en.wikipedia.org/wiki/Doris_Lessing
Doris Leuthard	http://en.wikipedia.org/wiki/Doris_Leuthard
Doris Roberts	http://en.wikipedia.org/wiki/Doris_Roberts
Doro Bush	http://en.wikipedia.org/wiki/Doro_Bush
Dorothea Dix	http://en.wikipedia.org/wiki/Dorothea_Dix
Dorothea Jordan	http://en.wikipedia.org/wiki/Dorothea_Jordan
Dorothea Lange	http://en.wikipedia.org/wiki/Dorothea_Lange
Dorothea Puente	http://en.wikipedia.org/wiki/Dorothea_Puente
Dorothy Allison	http://en.wikipedia.org/wiki/Dorothy_Allison
Dorothy Arzner	http://en.wikipedia.org/wiki/Dorothy_Arzner
Dorothy Canfield Fisher	http://en.wikipedia.org/wiki/Dorothy_Canfield_Fisher
Dorothy Crowfoot Hodgkin	http://en.wikipedia.org/wiki/Dorothy_Crowfoot_Hodgkin
Dorothy Dandridge	http://en.wikipedia.org/wiki/Dorothy_Dandridge
Dorothy Day	http://en.wikipedia.org/wiki/Dorothy_Day
Dorothy Denning	http://en.wikipedia.org/wiki/Dorothy_Denning
Dorothy Hamill	http://en.wikipedia.org/wiki/Dorothy_Hamill
Dorothy Kilgallen	http://en.wikipedia.org/wiki/Dorothy_Kilgallen
Dorothy L. Sayers	http://en.wikipedia.org/wiki/Dorothy_L._Sayers
Dorothy Lamour	http://en.wikipedia.org/wiki/Dorothy_Lamour
Dorothy Malone	http://en.wikipedia.org/wiki/Dorothy_Malone
Dorothy McGuire	http://en.wikipedia.org/wiki/Dorothy_McGuire
Dorothy Parker	http://en.wikipedia.org/wiki/Dorothy_Parker
Dorothy Richardson	http://en.wikipedia.org/wiki/Dorothy_Richardson
Dorothy Stickney	http://en.wikipedia.org/wiki/Dorothy_Stickney
Dorothy Stratten	http://en.wikipedia.org/wiki/Dorothy_Stratten
Dorothy Thompson	http://en.wikipedia.org/wiki/Dorothy_Thompson
Dorothy Tutin	http://en.wikipedia.org/wiki/Dorothy_Tutin
Dorothy West	http://en.wikipedia.org/wiki/Dorothy_West
Dorsey Burnette	http://en.wikipedia.org/wiki/Dorsey_Burnette
Dose One	http://en.wikipedia.org/wiki/Dose_One
Doug Barnard, Jr.	http://en.wikipedia.org/wiki/Doug_Barnard%2C_Jr.
Doug Bereuter	http://en.wikipedia.org/wiki/Doug_Bereuter
Doug Bereuter	http://en.wikipedia.org/wiki/Doug_Bereuter
Doug Coe	http://en.wikipedia.org/wiki/Doug_Coe
Doug E. Fresh	http://en.wikipedia.org/wiki/Doug_E._Fresh
Doug Engelbart	http://en.wikipedia.org/wiki/Doug_Engelbart
Doug Flutie	http://en.wikipedia.org/wiki/Doug_Flutie
Doug Henning	http://en.wikipedia.org/wiki/Doug_Henning
Doug Hutchison	http://en.wikipedia.org/wiki/Doug_Hutchison
Doug Lamborn	http://en.wikipedia.org/wiki/Doug_Lamborn
Doug McClure	http://en.wikipedia.org/wiki/Doug_McClure
Doug Ose	http://en.wikipedia.org/wiki/Doug_Ose
Doug Sahm	http://en.wikipedia.org/wiki/Doug_Sahm
Doug Savant	http://en.wikipedia.org/wiki/Doug_Savant
Doug Walgren	http://en.wikipedia.org/wiki/Doug_Walgren
Douglas Adams	http://en.wikipedia.org/wiki/Douglas_Adams
Douglas Alexander	http://en.wikipedia.org/wiki/Douglas_Alexander
Douglas Applegate	http://en.wikipedia.org/wiki/Douglas_Applegate
Douglas Carswell	http://en.wikipedia.org/wiki/Douglas_Carswell
Douglas Coupland	http://en.wikipedia.org/wiki/Douglas_Coupland
Douglas D. Osheroff	http://en.wikipedia.org/wiki/Douglas_D._Osheroff
Douglas Fairbanks, Jr.	http://en.wikipedia.org/wiki/Douglas_Fairbanks%2C_Jr.
Douglas Fairbanks, Sr.	http://en.wikipedia.org/wiki/Douglas_Fairbanks%2C_Sr.
Douglas Feith	http://en.wikipedia.org/wiki/Douglas_Feith
Douglas Fowley	http://en.wikipedia.org/wiki/Douglas_Fowley
Douglas H. Bosco	http://en.wikipedia.org/wiki/Douglas_H._Bosco
Douglas Hofstadter	http://en.wikipedia.org/wiki/Douglas_Hofstadter
Douglas Kennedy	http://en.wikipedia.org/wiki/Douglas_Kennedy_(actor)
Douglas Lowenstein	http://en.wikipedia.org/wiki/Douglas_Lowenstein
Douglas MacArthur	http://en.wikipedia.org/wiki/Douglas_MacArthur
Douglas McKay	http://en.wikipedia.org/wiki/Douglas_McKay
Douglas Rushkoff	http://en.wikipedia.org/wiki/Douglas_Rushkoff
Douglas Sirk	http://en.wikipedia.org/wiki/Douglas_Sirk
Douglas Stewart	http://en.wikipedia.org/wiki/Douglas_Stewart
Douglas Stuart Moore	http://en.wikipedia.org/wiki/Douglas_Stuart_Moore
Douglas Trumbull	http://en.wikipedia.org/wiki/Douglas_Trumbull
Douglas W. Kmiec	http://en.wikipedia.org/wiki/Douglas_W._Kmiec
Douglas Wilson	http://en.wikipedia.org/wiki/Douglas_Wilson_(interior_designer)
Douglas Woolf	http://en.wikipedia.org/wiki/Douglas_Woolf
Dougray Scott	http://en.wikipedia.org/wiki/Dougray_Scott
Dov Charney	http://en.wikipedia.org/wiki/Dov_Charney
Downtown Julie Brown	http://en.wikipedia.org/wiki/Downtown_Julie_Brown
Doyle McManus	http://en.wikipedia.org/wiki/Doyle_McManus
Dr. Dean Edell	http://en.wikipedia.org/wiki/Dr._Dean_Edell
Dr. Demento	http://en.wikipedia.org/wiki/Dr._Demento
Dr. Dre	http://en.wikipedia.org/wiki/Dr._Dre
Dr. Gene Scott	http://en.wikipedia.org/wiki/Dr._Gene_Scott
Dr. Michael Baden	http://en.wikipedia.org/wiki/Dr._Michael_Baden
Dr. Neal Barnard	http://en.wikipedia.org/wiki/Dr._Neal_Barnard
Dr. Ralph Stanley	http://en.wikipedia.org/wiki/Dr._Ralph_Stanley
Dr. Seuss	http://en.wikipedia.org/wiki/Dr._Seuss
Dragan Cavic	http://en.wikipedia.org/wiki/Dragan_Cavic
Drake Bell	http://en.wikipedia.org/wiki/Drake_Bell
Drea de Matteo	http://en.wikipedia.org/wiki/Drea_de_Matteo
Drew Barrymore	http://en.wikipedia.org/wiki/Drew_Barrymore
Drew Bledsoe	http://en.wikipedia.org/wiki/Drew_Bledsoe
Drew Brees	http://en.wikipedia.org/wiki/Drew_Brees
Drew Carey	http://en.wikipedia.org/wiki/Drew_Carey
Drew Curtis	http://en.wikipedia.org/wiki/Drew_Curtis
Drew Daniel	http://en.wikipedia.org/wiki/Andrew_Daniel
Drew Fuller	http://en.wikipedia.org/wiki/Drew_Fuller
Drew Lewis	http://en.wikipedia.org/wiki/Drew_Lewis
Drew Pearson	http://en.wikipedia.org/wiki/Drew_Pearson_(journalist)
Driss Jettou	http://en.wikipedia.org/wiki/Driss_Jettou
Duane Allman	http://en.wikipedia.org/wiki/Duane_Allman
Duane Denison	http://en.wikipedia.org/wiki/Duane_Denison
Duane Eddy	http://en.wikipedia.org/wiki/Duane_Eddy
Duane Jones	http://en.wikipedia.org/wiki/Duane_Jones
Duane Martin	http://en.wikipedia.org/wiki/Duane_Martin
DuBose Heyward	http://en.wikipedia.org/wiki/DuBose_Heyward
Duccio di Buoninsegna	http://en.wikipedia.org/wiki/Duccio_di_Buoninsegna
Dudley Fitts	http://en.wikipedia.org/wiki/Dudley_Fitts
Dudley Moore	http://en.wikipedia.org/wiki/Dudley_Moore
Dudley R. Herschbach	http://en.wikipedia.org/wiki/Dudley_R._Herschbach
Duff Green	http://en.wikipedia.org/wiki/Duff_Green
Duff McKagan	http://en.wikipedia.org/wiki/Duff_McKagan
Duke Cunningham	http://en.wikipedia.org/wiki/Duke_Cunningham
Duke Ellington	http://en.wikipedia.org/wiki/Duke_Ellington
Duke Snider	http://en.wikipedia.org/wiki/Duke_Snider
Dul� Hill	http://en.wikipedia.org/wiki/Dul%C3%A9_Hill
Dumas Malone	http://en.wikipedia.org/wiki/Dumas_Malone
Duncan D. Hunter	http://en.wikipedia.org/wiki/Duncan_D._Hunter
Duncan Hames	http://en.wikipedia.org/wiki/Duncan_Hames
Duncan Hunter	http://en.wikipedia.org/wiki/Duncan_Hunter
Duncan I	http://en.wikipedia.org/wiki/Duncan_I
Duncan II	http://en.wikipedia.org/wiki/Duncan_II
Duncan Sheik	http://en.wikipedia.org/wiki/Duncan_Sheik
Dustin Diamond	http://en.wikipedia.org/wiki/Dustin_Diamond
Dustin Hoffman	http://en.wikipedia.org/wiki/Dustin_Hoffman
Dusty Springfield	http://en.wikipedia.org/wiki/Dusty_Springfield
Dutch Ruppersberger	http://en.wikipedia.org/wiki/Dusty_Springfield
Dwayne Andreas	http://en.wikipedia.org/wiki/Dwayne_Andreas
Dwayne Goettel	http://en.wikipedia.org/wiki/Dwayne_Goettel
Dwayne Hickman	http://en.wikipedia.org/wiki/Dwayne_Hickman
Dweezil Zappa	http://en.wikipedia.org/wiki/Dweezil_Zappa
Dwight D. Eisenhower	http://en.wikipedia.org/wiki/Dwight_D._Eisenhower
Dwight Gooden	http://en.wikipedia.org/wiki/Dwight_Gooden
Dwight Macdonald	http://en.wikipedia.org/wiki/Dwight_Macdonald
Dwight Schultz	http://en.wikipedia.org/wiki/Dwight_Schultz
Dwight Yoakam	http://en.wikipedia.org/wiki/Dwight_Yoakam
Dwight Yoakam	http://en.wikipedia.org/wiki/Dwight_Yoakam
Dwyane Wade	http://en.wikipedia.org/wiki/Dwyane_Wade
Dyan Cannon	http://en.wikipedia.org/wiki/Dyan_Cannon
Dylan Klebold	http://en.wikipedia.org/wiki/Dylan_Klebold
Dylan McDermott	http://en.wikipedia.org/wiki/Dylan_McDermott
Dylan Moran	http://en.wikipedia.org/wiki/Dylan_Moran
Dylan Sprouse	http://en.wikipedia.org/wiki/Dylan_Sprouse
Dylan Thomas	http://en.wikipedia.org/wiki/Dylan_Thomas
Dylan Walsh	http://en.wikipedia.org/wiki/Dylan_Walsh
Dzhokhar Dudayev	http://en.wikipedia.org/wiki/Dzhokhar_Dudayev
E. Annie Proulx	http://en.wikipedia.org/wiki/E._Annie_Proulx
E. B. White	http://en.wikipedia.org/wiki/E._B._White
E. Clay Shaw	http://en.wikipedia.org/wiki/E._Clay_Shaw
E. Clay Shaw, Jr.	http://en.wikipedia.org/wiki/E._Clay_Shaw%2C_Jr.
E. E. "Doc" Smith	http://en.wikipedia.org/wiki/E._E._%22Doc%22_Smith
e. e. cummings	http://en.wikipedia.org/wiki/e._e._cummings
E. Franklin Frazier	http://en.wikipedia.org/wiki/E._Franklin_Frazier
E. G. Marshall	http://en.wikipedia.org/wiki/E._G._Marshall
E. H. Gombrich	http://en.wikipedia.org/wiki/E._H._Gombrich
E. Howard Hunt	http://en.wikipedia.org/wiki/E._Howard_Hunt
E. J. Dionne	http://en.wikipedia.org/wiki/E._Howard_Hunt
E. J. Pratt	http://en.wikipedia.org/wiki/E._J._Pratt
E. L. Doctorow	http://en.wikipedia.org/wiki/E._L._Doctorow
E. L. Godkin	http://en.wikipedia.org/wiki/E._L._Godkin
E. M. Forster	http://en.wikipedia.org/wiki/E._M._Forster
E. M. Purcell	http://en.wikipedia.org/wiki/E._M._Purcell
E. Nesbit	http://en.wikipedia.org/wiki/E._Nesbit
E. P. Thompson	http://en.wikipedia.org/wiki/E._P._Thompson
E. Parry Thomas	http://en.wikipedia.org/wiki/E._Parry_Thomas
E. R. Braithwaite	http://en.wikipedia.org/wiki/E._R._Braithwaite
E. Stanley O'Neal	http://en.wikipedia.org/wiki/E._Stanley_O%27Neal
E. T. A. Hoffmann	http://en.wikipedia.org/wiki/E._T._A._Hoffmann
E. V. Knox	http://en.wikipedia.org/wiki/E._V._Knox
E. Z. C. Judson	http://en.wikipedia.org/wiki/E._Z._C._Judson
Eadweard Muybridge	http://en.wikipedia.org/wiki/Eadweard_Muybridge
Eagle-Eye Cherry	http://en.wikipedia.org/wiki/Eagle-Eye_Cherry
Eamon de Valera	http://en.wikipedia.org/wiki/Eamon_de_Valera
Earl Anthony	http://en.wikipedia.org/wiki/Earl_Anthony
Earl Blumenauer	http://en.wikipedia.org/wiki/Earl_Blumenauer
Earl Boen	http://en.wikipedia.org/wiki/Earl_Boen
Earl Butz	http://en.wikipedia.org/wiki/Earl_Butz
Earl Campbell	http://en.wikipedia.org/wiki/Earl_Campbell
Earl Hilliard	http://en.wikipedia.org/wiki/Earl_Hilliard
Earl Hindman	http://en.wikipedia.org/wiki/Earl_Hindman
Earl Holliman	http://en.wikipedia.org/wiki/Earl_Holliman
Earl Hutto	http://en.wikipedia.org/wiki/Earl_Hutto
Earl Pomeroy	http://en.wikipedia.org/wiki/Earl_Pomeroy
Earl Scruggs	http://en.wikipedia.org/wiki/Earl_Scruggs
Earl Warren	http://en.wikipedia.org/wiki/Earl_Warren
Earle Birney	http://en.wikipedia.org/wiki/Earle_Birney
Earle Brown	http://en.wikipedia.org/wiki/Earle_Brown
Eartha Kitt	http://en.wikipedia.org/wiki/Eartha_Kitt
Eavan Boland	http://en.wikipedia.org/wiki/Eavan_Boland
Eberhard Weber	http://en.wikipedia.org/wiki/Eberhard_Weber
Eckhard Pfeiffer	http://en.wikipedia.org/wiki/Eckhard_Pfeiffer
Ed Altman	http://en.wikipedia.org/wiki/Edward_Altman
Ed Ames	http://en.wikipedia.org/wiki/Ed_Ames
Ed Asner	http://en.wikipedia.org/wiki/Ed_Asner
Ed Balls	http://en.wikipedia.org/wiki/Ed_Balls
Ed Begley, Jr.	http://en.wikipedia.org/wiki/Ed_Begley%2C_Jr.
Ed Begley, Sr.	http://en.wikipedia.org/wiki/Ed_Begley%2C_Sr.
Ed Bethune	http://en.wikipedia.org/wiki/Ed_Bethune
Ed Bradley	http://en.wikipedia.org/wiki/Ed_Bradley
Ed Buckham	http://en.wikipedia.org/wiki/Ed_Buckham
Ed Bullins	http://en.wikipedia.org/wiki/Ed_Bullins
Ed Case	http://en.wikipedia.org/wiki/Ed_Case
Ed Felten	http://en.wikipedia.org/wiki/Ed_Felten
Ed Flanders	http://en.wikipedia.org/wiki/Ed_Flanders
Ed Gein	http://en.wikipedia.org/wiki/Ed_Gein
Ed Gillespie	http://en.wikipedia.org/wiki/Ed_Gillespie
Ed Guthman	http://en.wikipedia.org/wiki/Ed_Guthman
Ed Harris	http://en.wikipedia.org/wiki/Ed_Harris
Ed Helms	http://en.wikipedia.org/wiki/Ed_Helms
Ed Jenkins	http://en.wikipedia.org/wiki/Ed_Jenkins_(politician)
Ed Jones	http://en.wikipedia.org/wiki/Ed_Jones_(U.S._politician)
Ed Kemper	http://en.wikipedia.org/wiki/Ed_Kemper
Ed Koch	http://en.wikipedia.org/wiki/Ed_Koch
Ed Marinaro	http://en.wikipedia.org/wiki/Ed_Marinaro
Ed Markey	http://en.wikipedia.org/wiki/Ed_Markey
Ed McMahon	http://en.wikipedia.org/wiki/Ed_McMahon
Ed Meese	http://en.wikipedia.org/wiki/Ed_Meese
Ed Miliband	http://en.wikipedia.org/wiki/Ed_Miliband
Ed Muskie	http://en.wikipedia.org/wiki/Ed_Muskie
Ed O'Brien	http://en.wikipedia.org/wiki/Ed_O%27Brien
Ed O'Neill	http://en.wikipedia.org/wiki/Ed_O%27Neill
Ed Pastor	http://en.wikipedia.org/wiki/Ed_Pastor
Ed Perlmutter	http://en.wikipedia.org/wiki/Ed_Perlmutter
Ed Rendell	http://en.wikipedia.org/wiki/Ed_Rendell
Ed Rendell	http://en.wikipedia.org/wiki/Ed_Rendell
Ed Rollins	http://en.wikipedia.org/wiki/Ed_Rollins
Ed Royce	http://en.wikipedia.org/wiki/Ed_Royce
Ed Simons	http://en.wikipedia.org/wiki/Ed_Simons
Ed Sullivan	http://en.wikipedia.org/wiki/Ed_Sullivan
Ed Templeton	http://en.wikipedia.org/wiki/Ed_Templeton
Ed Townsend	http://en.wikipedia.org/wiki/Ed_Townsend
Ed Whitacre, Jr.	http://en.wikipedia.org/wiki/Ed_Whitacre%2C_Jr.
Ed White	http://en.wikipedia.org/wiki/Edward_Higgins_White
Ed Whitfield	http://en.wikipedia.org/wiki/Ed_Whitfield
Ed Wood	http://en.wikipedia.org/wiki/Ed_Wood
Ed Wynn	http://en.wikipedia.org/wiki/Ed_Wynn
Ed Zander	http://en.wikipedia.org/wiki/Ed_Zander
Ed Zschau	http://en.wikipedia.org/wiki/Ed_Zschau
Eddie Albert	http://en.wikipedia.org/wiki/Eddie_Albert
Eddie Antar	http://en.wikipedia.org/wiki/Eddie_Antar
Eddie Arcaro	http://en.wikipedia.org/wiki/Eddie_Arcaro
Eddie Bernice Johnson	http://en.wikipedia.org/wiki/Eddie_Bernice_Johnson
Eddie Bracken	http://en.wikipedia.org/wiki/Eddie_Bracken
Eddie Campbell	http://en.wikipedia.org/wiki/Eddie_Campbell
Eddie Cantor	http://en.wikipedia.org/wiki/Eddie_Cantor
Eddie Cibrian	http://en.wikipedia.org/wiki/Eddie_Cibrian
Eddie Cochran	http://en.wikipedia.org/wiki/Eddie_Cochran
Eddie Collins	http://en.wikipedia.org/wiki/Eddie_Collins
Eddie DeBartolo, Jr.	http://en.wikipedia.org/wiki/Eddie_DeBartolo%2C_Jr.
Eddie Deezen	http://en.wikipedia.org/wiki/Eddie_Deezen
Eddie Fenech Adami	http://en.wikipedia.org/wiki/Eddie_Fenech_Adami
Eddie Fisher	http://en.wikipedia.org/wiki/Eddie_Fisher_(singer)
Eddie Floyd	http://en.wikipedia.org/wiki/Eddie_Floyd
Eddie Fontaine	http://en.wikipedia.org/wiki/Eddie_Fontaine
Eddie Furlong	http://en.wikipedia.org/wiki/Eddie_Furlong
Eddie Griffin	http://en.wikipedia.org/wiki/Eddie_Griffin
Eddie Guerrero	http://en.wikipedia.org/wiki/Eddie_Guerrero
Eddie Holland	http://en.wikipedia.org/wiki/Eddie_Holland
Eddie Izzard	http://en.wikipedia.org/wiki/Eddie_Izzard
Eddie Kendricks	http://en.wikipedia.org/wiki/Eddie_Kendricks
Eddie Mathews	http://en.wikipedia.org/wiki/Eddie_Mathews
Eddie Money	http://en.wikipedia.org/wiki/Eddie_Money
Eddie Murphy	http://en.wikipedia.org/wiki/Eddie_Murphy
Eddie Murray	http://en.wikipedia.org/wiki/Eddie_Murray
Eddie Quillan	http://en.wikipedia.org/wiki/Eddie_Quillan
Eddie Rabbitt	http://en.wikipedia.org/wiki/Eddie_Rabbitt
Eddie Rickenbacker	http://en.wikipedia.org/wiki/Eddie_Rickenbacker
Eddie Slovik	http://en.wikipedia.org/wiki/Eddie_Slovik
Eddie Van Halen	http://en.wikipedia.org/wiki/Eddie_Van_Halen
Eddie Vedder	http://en.wikipedia.org/wiki/Eddie_Vedder
Eddy Arnold	http://en.wikipedia.org/wiki/Eddy_Arnold
Eddy Grant	http://en.wikipedia.org/wiki/Eddy_Grant
Ede Szigligeti	http://en.wikipedia.org/wiki/Ede_Szigligeti
Edem Kodjo	http://en.wikipedia.org/wiki/Edem_Kodjo
Edgar Allan Poe	http://en.wikipedia.org/wiki/Edgar_Allan_Poe
Edgar Atheling	http://en.wikipedia.org/wiki/Edgar_Atheling
Edgar Bergen	http://en.wikipedia.org/wiki/Edgar_Bergen
Edgar Bowers	http://en.wikipedia.org/wiki/Edgar_Bowers
Edgar Bronfman, Jr.	http://en.wikipedia.org/wiki/Edgar_Bronfman%2C_Jr.
Edgar Bronfman, Sr.	http://en.wikipedia.org/wiki/Edgar_Bronfman%2C_Sr.
Edgar Buchanan	http://en.wikipedia.org/wiki/Edgar_Buchanan
Edgar Cayce	http://en.wikipedia.org/wiki/Edgar_Cayce
Edgar Degas	http://en.wikipedia.org/wiki/Edgar_Degas
Edgar Guest	http://en.wikipedia.org/wiki/Edgar_Guest
Edgar Kennedy	http://en.wikipedia.org/wiki/Edgar_Kennedy
Edgar Lee Masters	http://en.wikipedia.org/wiki/Edgar_Lee_Masters
Edgar Ray Killen	http://en.wikipedia.org/wiki/Edgar_Ray_Killen
Edgar Rice Burroughs	http://en.wikipedia.org/wiki/Edgar_Rice_Burroughs
Edgar Wallace	http://en.wikipedia.org/wiki/Edgar_Wallace
Edgar Winter	http://en.wikipedia.org/wiki/Edgar_Winter
Edgard Var�se	http://en.wikipedia.org/wiki/Edgard_Var%C3%A8se
Edie Adams	http://en.wikipedia.org/wiki/Edie_Adams
Edie Brickell	http://en.wikipedia.org/wiki/Edie_Brickell
Edie Falco	http://en.wikipedia.org/wiki/Edie_Falco
Edie McClurg	http://en.wikipedia.org/wiki/Edie_McClurg
Edith Cresson	http://en.wikipedia.org/wiki/Edith_Cresson
Edith Evans	http://en.wikipedia.org/wiki/Edith_Evans
Edith Hamilton	http://en.wikipedia.org/wiki/Edith_Hamilton
Edith Jones	http://en.wikipedia.org/wiki/Edith_Jones
Edith Piaf	http://en.wikipedia.org/wiki/Edith_Piaf
Edith Sitwell	http://en.wikipedia.org/wiki/Edith_Sitwell
Edith Wharton	http://en.wikipedia.org/wiki/Edith_Wharton
Edme Mariotte	http://en.wikipedia.org/wiki/Edme_Mariotte
Edmond Fr�my	http://en.wikipedia.org/wiki/Edmond_Fr%C3%A9my
Edmond Hoyle	http://en.wikipedia.org/wiki/Edmond_Hoyle
Edmond Malone	http://en.wikipedia.org/wiki/Edmond_Malone
Edmond O'Brien	http://en.wikipedia.org/wiki/Edmond_O%27Brien
Edmond Rostand	http://en.wikipedia.org/wiki/Edmond_Rostand
Edmund Allenby	http://en.wikipedia.org/wiki/Edmund_Allenby
Edmund Andros	http://en.wikipedia.org/wiki/Edmund_Andros
Edmund Beecher Wilson	http://en.wikipedia.org/wiki/Edmund_Beecher_Wilson
Edmund Blunden	http://en.wikipedia.org/wiki/Edmund_Blunden
Edmund Bolton	http://en.wikipedia.org/wiki/Edmund_Bolton
Edmund Burke	http://en.wikipedia.org/wiki/Edmund_Burke
Edmund Cartwright	http://en.wikipedia.org/wiki/Edmund_Cartwright
Edmund Castell	http://en.wikipedia.org/wiki/Edmund_Castell
Edmund Curll	http://en.wikipedia.org/wiki/Edmund_Curll
Edmund Dulac	http://en.wikipedia.org/wiki/Edmund_Dulac
Edmund Goulding	http://en.wikipedia.org/wiki/Edmund_Goulding
Edmund Gwenn	http://en.wikipedia.org/wiki/Edmund_Gwenn
Edmund Halley	http://en.wikipedia.org/wiki/Edmund_Halley
Edmund Hillary	http://en.wikipedia.org/wiki/Edmund_Hillary
Edmund Ho	http://en.wikipedia.org/wiki/Edmund_Ho
Edmund Husserl	http://en.wikipedia.org/wiki/Edmund_Husserl
Edmund Kean	http://en.wikipedia.org/wiki/Edmund_Kean
Edmund Kirby Smith	http://en.wikipedia.org/wiki/Edmund_Kirby_Smith
Edmund Ludlow	http://en.wikipedia.org/wiki/Edmund_Ludlow
Edmund Randolph	http://en.wikipedia.org/wiki/Edmund_Randolph
Edmund Spenser	http://en.wikipedia.org/wiki/Edmund_Spenser
Edmund Waller	http://en.wikipedia.org/wiki/Edmund_Waller
Edmund White	http://en.wikipedia.org/wiki/Edmund_White
Edmund Wilson	http://en.wikipedia.org/wiki/Edmund_Wilson
Edna Best	http://en.wikipedia.org/wiki/Edna_Best
Edna Ferber	http://en.wikipedia.org/wiki/Edna_Ferber
Edna O'Brien	http://en.wikipedia.org/wiki/Edna_O%27Brien
Edna St. Vincent Millay	http://en.wikipedia.org/wiki/Edna_St._Vincent_Millay
Edolphus Towns	http://en.wikipedia.org/wiki/Edolphus_Towns
Edolphus Towns	http://en.wikipedia.org/wiki/Edolphus_Towns
�douard Balladur	http://en.wikipedia.org/wiki/%C9douard_Balladur
�douard Daladier	http://en.wikipedia.org/wiki/%C9douard_Daladier
�douard Glissant	http://en.wikipedia.org/wiki/%C9douard_Glissant
Edouard Manet	http://en.wikipedia.org/wiki/Edouard_Manet
Edsel Ford	http://en.wikipedia.org/wiki/Edsel_Ford
Edsger Dijkstra	http://en.wikipedia.org/wiki/Edsger_Dijkstra
Eduard Benes	http://en.wikipedia.org/wiki/Eduard_Benes
Eduard Buchner	http://en.wikipedia.org/wiki/Eduard_Buchner
Eduard Kokoyty	http://en.wikipedia.org/wiki/Eduard_Kokoyty
Eduard Shevardnadze	http://en.wikipedia.org/wiki/Eduard_Shevardnadze
Eduard Suess	http://en.wikipedia.org/wiki/Eduard_Suess
Eduard von Hartmann	http://en.wikipedia.org/wiki/Eduard_von_Hartmann
Eduardo Paolozzi	http://en.wikipedia.org/wiki/Eduardo_Paolozzi
Eduardo Rodriguez	http://en.wikipedia.org/wiki/Eduardo_Rodríguez
Eduardo Verastegui	http://en.wikipedia.org/wiki/Eduardo_Verastegui
Edvard Grieg	http://en.wikipedia.org/wiki/Edvard_Grieg
Edvard Munch	http://en.wikipedia.org/wiki/Edvard_Munch
Edvard Westermarck	http://en.wikipedia.org/wiki/Edvard_Westermarck
Edward Abbey	http://en.wikipedia.org/wiki/Edward_Abbey
Edward Addison	http://en.wikipedia.org/wiki/Edward_Addison
Edward Albee	http://en.wikipedia.org/wiki/Edward_Albee
Edward Albert	http://en.wikipedia.org/wiki/Edward_Albert
Edward Arnold	http://en.wikipedia.org/wiki/Edward_Arnold_(actor)
Edward Artemiev	http://en.wikipedia.org/wiki/Edward_Artemiev
Edward B. Lewis	http://en.wikipedia.org/wiki/Edward_B._Lewis
Edward Bernays	http://en.wikipedia.org/wiki/Edward_Bernays
Edward Binns	http://en.wikipedia.org/wiki/Edward_Binns
Edward Bok	http://en.wikipedia.org/wiki/Edward_Bok
Edward Bond	http://en.wikipedia.org/wiki/Edward_Bond
Edward Boscawen	http://en.wikipedia.org/wiki/Edward_Boscawen
Edward Braddock	http://en.wikipedia.org/wiki/Edward_Braddock
Edward Bunker	http://en.wikipedia.org/wiki/Edward_Bunker
Edward Burne-Jones	http://en.wikipedia.org/wiki/Edward_Burne-Jones
Edward Burns	http://en.wikipedia.org/wiki/Edward_Burns
Edward Channing	http://en.wikipedia.org/wiki/Edward_Channing
Edward Charles Pickering	http://en.wikipedia.org/wiki/Edward_Charles_Pickering
Edward Cox	http://en.wikipedia.org/wiki/Edward_F._Cox
Edward Dahlberg	http://en.wikipedia.org/wiki/Edward_Dahlberg
Edward Davey	http://en.wikipedia.org/wiki/Edward_Davey
Edward Dmytryk	http://en.wikipedia.org/wiki/Edward_Dmytryk
Edward Drinker Cope	http://en.wikipedia.org/wiki/Edward_Drinker_Cope
Edward Eggleston	http://en.wikipedia.org/wiki/Edward_Eggleston
Edward Elgar	http://en.wikipedia.org/wiki/Edward_Elgar
Edward Evans-Pritchard	http://en.wikipedia.org/wiki/Edward_Evans-Pritchard
Edward Everett Hale	http://en.wikipedia.org/wiki/Edward_Everett_Hale
Edward Everett Horton	http://en.wikipedia.org/wiki/Edward_Everett_Horton
Edward F. Feighan	http://en.wikipedia.org/wiki/Edward_F._Feighan
Edward Forbes	http://en.wikipedia.org/wiki/Edward_Forbes
Edward Fox	http://en.wikipedia.org/wiki/Edward_Fox_(actor)
Edward Furlong	http://en.wikipedia.org/wiki/Edward_Furlong
Edward G. Robinson	http://en.wikipedia.org/wiki/Edward_G._Robinson
Edward Garnier	http://en.wikipedia.org/wiki/Edward_Garnier
Edward George Bulwer-Lytton	http://en.wikipedia.org/wiki/Edward_George_Bulwer-Lytton
Edward Gibbon	http://en.wikipedia.org/wiki/Edward_Gibbon
Edward Gibbon Wakefield	http://en.wikipedia.org/wiki/Edward_Gibbon_Wakefield
Edward Gorey	http://en.wikipedia.org/wiki/Edward_Gorey
Edward Hall	http://en.wikipedia.org/wiki/Edward_Hall
Edward Hawke	http://en.wikipedia.org/wiki/Edward_Hawke
Edward Heath	http://en.wikipedia.org/wiki/Edward_Heath
Edward Herrmann	http://en.wikipedia.org/wiki/Edward_Herrmann
Edward Hibbert	http://en.wikipedia.org/wiki/Edward_Hibbert
Edward Hoagland	http://en.wikipedia.org/wiki/Edward_Hoagland
Edward Hopper	http://en.wikipedia.org/wiki/Edward_Hopper
Edward Horsman	http://en.wikipedia.org/wiki/Edward_Horsman
Edward Irving	http://en.wikipedia.org/wiki/Edward_Irving
Edward J. Markey	http://en.wikipedia.org/wiki/Edward_J._Markey
Edward J. Piszek	http://en.wikipedia.org/wiki/Edward_Piszek
Edward James Olmos	http://en.wikipedia.org/wiki/Edward_James_Olmos
Edward Jenner	http://en.wikipedia.org/wiki/Edward_Jenner
Edward Ka-Spel	http://en.wikipedia.org/wiki/Edward_Ka-Spel
Edward L. Schrock	http://en.wikipedia.org/wiki/Edward_L._Schrock
Edward Lear	http://en.wikipedia.org/wiki/Edward_Lear
Edward Leigh	http://en.wikipedia.org/wiki/Edward_Leigh
Edward Livingston	http://en.wikipedia.org/wiki/Edward_Livingston
Edward Lowassa	http://en.wikipedia.org/wiki/Edward_Lowassa
Edward M. House	http://en.wikipedia.org/wiki/Edward_M._House
Edward M. Kennedy	http://en.wikipedia.org/wiki/Edward_M._Kennedy
Edward MacDowell	http://en.wikipedia.org/wiki/Edward_MacDowell
Edward Madigan	http://en.wikipedia.org/wiki/Edward_Madigan
Edward Miliband	http://en.wikipedia.org/wiki/Edward_Miliband
Edward Mulhare	http://en.wikipedia.org/wiki/Edward_Mulhare
Edward Natapei	http://en.wikipedia.org/wiki/Edward_Natapei
Edward Norton	http://en.wikipedia.org/wiki/Edward_Norton
Edward Noyes Westcott	http://en.wikipedia.org/wiki/Edward_Noyes_Westcott
Edward O. Wilson	http://en.wikipedia.org/wiki/Edward_O._Wilson
Edward P. Boland	http://en.wikipedia.org/wiki/Edward_P._Boland
Edward P. Jones	http://en.wikipedia.org/wiki/Edward_P._Jones
Edward R. Murrow	http://en.wikipedia.org/wiki/Edward_R._Murrow
Edward R. Roybal	http://en.wikipedia.org/wiki/Edward_R._Roybal
Edward R. Roybal	http://en.wikipedia.org/wiki/Edward_R._Roybal
Edward Ruscha	http://en.wikipedia.org/wiki/Edward_Ruscha
Edward Said	http://en.wikipedia.org/wiki/Edward_Said
Edward Sapir	http://en.wikipedia.org/wiki/Edward_Sapir
Edward Schillebeeckx	http://en.wikipedia.org/wiki/Edward_Schillebeeckx
Edward Steichen	http://en.wikipedia.org/wiki/Edward_Steichen
Edward Stettinius, Jr.	http://en.wikipedia.org/wiki/Edward_Stettinius%2C_Jr.
Edward Teller	http://en.wikipedia.org/wiki/Edward_Teller
Edward the Black Prince	http://en.wikipedia.org/wiki/Edward_the_Black_Prince
Edward the Confessor	http://en.wikipedia.org/wiki/Edward_the_Confessor
Edward the Martyr	http://en.wikipedia.org/wiki/Edward_the_Martyr
Edward Timpson	http://en.wikipedia.org/wiki/Edward_Timpson
Edward Tufte	http://en.wikipedia.org/wiki/Edward_Tufte
Edward Tylor	http://en.wikipedia.org/wiki/Edward_Tylor
Edward Vaizey	http://en.wikipedia.org/wiki/Edward_Vaizey
Edward Victor Appleton	http://en.wikipedia.org/wiki/Edward_Victor_Appleton
Edward Villella	http://en.wikipedia.org/wiki/Edward_Villella
Edward Walker	http://en.wikipedia.org/wiki/Edward_S._Walker,_Jr.
Edward Whymper	http://en.wikipedia.org/wiki/Edward_Whymper
Edward Winslow	http://en.wikipedia.org/wiki/Edward_Winslow
Edward Woodward	http://en.wikipedia.org/wiki/Edward_Woodward
Edward Young	http://en.wikipedia.org/wiki/Edward_Young
Edward Zorinsky	http://en.wikipedia.org/wiki/Edward_Zorinsky
Edwidge Danticat	http://en.wikipedia.org/wiki/Edwidge_Danticat
Edwin Alonzo Boyd	http://en.wikipedia.org/wiki/Edwin_Alonzo_Boyd
Edwin Arlington Robinson	http://en.wikipedia.org/wiki/Edwin_Arlington_Robinson
Edwin Edwards	http://en.wikipedia.org/wiki/Edwin_Edwards
Edwin Feulner	http://en.wikipedia.org/wiki/Edwin_Feulner
Edwin Forrest	http://en.wikipedia.org/wiki/Edwin_Forrest
Edwin G. Boring	http://en.wikipedia.org/wiki/Edwin_G._Boring
Edwin H. Armstrong	http://en.wikipedia.org/wiki/Edwin_H._Armstrong
Edwin Hall	http://en.wikipedia.org/wiki/Edwin_Hall
Edwin Hubble	http://en.wikipedia.org/wiki/Edwin_Hubble
Edwin Lutyens	http://en.wikipedia.org/wiki/Edwin_Lutyens
Edwin M. McMillan	http://en.wikipedia.org/wiki/Edwin_M._McMillan
Edwin M. Stanton	http://en.wikipedia.org/wiki/Edwin_M._Stanton
Edwin Markham	http://en.wikipedia.org/wiki/Edwin_Markham
Edwin Moses	http://en.wikipedia.org/wiki/Edwin_Moses
Edwin Moses	http://en.wikipedia.org/wiki/Edwin_Moses
Edwin Newman	http://en.wikipedia.org/wiki/Edwin_Newman
Edwin O'Connor	http://en.wikipedia.org/wiki/Edwin_O%27Connor
Edwin Starr	http://en.wikipedia.org/wiki/Edwin_Starr
Edwin Vose Sumner	http://en.wikipedia.org/wiki/Edwin_Vose_Sumner
Eero Saarinen	http://en.wikipedia.org/wiki/Eero_Saarinen
Efraim Halevy	http://en.wikipedia.org/wiki/Efraim_Halevy
Efrem Zimbalist, Jr.	http://en.wikipedia.org/wiki/Efrem_Zimbalist%2C_Jr.
Egon Krenz	http://en.wikipedia.org/wiki/Egon_Krenz
Egon Schiele	http://en.wikipedia.org/wiki/Egon_Schiele
Ehud Barak	http://en.wikipedia.org/wiki/Ehud_Barak
Ehud Olmert	http://en.wikipedia.org/wiki/Ehud_Olmert
Ehud Olmert	http://en.wikipedia.org/wiki/Ehud_Olmert
Eileen Atkins	http://en.wikipedia.org/wiki/Eileen_Atkins
Eileen Brennan	http://en.wikipedia.org/wiki/Eileen_Brennan
Eileen Heckart	http://en.wikipedia.org/wiki/Eileen_Heckart
Eilidh Whiteford	http://en.wikipedia.org/wiki/Eilidh_Whiteford
Einar Orn	http://en.wikipedia.org/wiki/Einar_Orn
Eion Bailey	http://en.wikipedia.org/wiki/Eion_Bailey
Eisaku Sato	http://en.wikipedia.org/wiki/Eisaku_Sato
El DeBarge	http://en.wikipedia.org/wiki/El_DeBarge
El Greco	http://en.wikipedia.org/wiki/El_Greco
Elaine Chao	http://en.wikipedia.org/wiki/Elaine_Chao
Elaine Joyce	http://en.wikipedia.org/wiki/Elaine_Joyce
Elaine May	http://en.wikipedia.org/wiki/Elaine_May
Elaine Miles	http://en.wikipedia.org/wiki/Elaine_Miles
Elaine Showalter	http://en.wikipedia.org/wiki/Elaine_Showalter
Elaine Stritch	http://en.wikipedia.org/wiki/Elaine_Stritch
Elayne Boosler	http://en.wikipedia.org/wiki/Elayne_Boosler
Elbert Henry Gary	http://en.wikipedia.org/wiki/Elbert_Henry_Gary
Elbert Hubbard	http://en.wikipedia.org/wiki/Elbert_Hubbard
Elbridge Bryant	http://en.wikipedia.org/wiki/Elbridge_Bryant
Elbridge Gerry	http://en.wikipedia.org/wiki/Elbridge_Gerry
Elden Henson	http://en.wikipedia.org/wiki/Elden_Henson
Eldon Dedini	http://en.wikipedia.org/wiki/Eldon_Dedini
Eldon Rudd	http://en.wikipedia.org/wiki/Eldon_Rudd
Eldridge Cleaver	http://en.wikipedia.org/wiki/Eldridge_Cleaver
Eleanor H. Porter	http://en.wikipedia.org/wiki/Eleanor_H._Porter
Eleanor Holmes Norton	http://en.wikipedia.org/wiki/Eleanor_Holmes_Norton
Eleanor Laing	http://en.wikipedia.org/wiki/Eleanor_Laing
Eleanor of Aquitaine	http://en.wikipedia.org/wiki/Eleanor_of_Aquitaine
Eleanor Parker	http://en.wikipedia.org/wiki/Eleanor_Parker
Eleanor Powell	http://en.wikipedia.org/wiki/Eleanor_Powell
Eleanor Roosevelt	http://en.wikipedia.org/wiki/Eleanor_Roosevelt
Eleanora Duse	http://en.wikipedia.org/wiki/Eleanora_Duse
Elena Poniatowska	http://en.wikipedia.org/wiki/Elena_Poniatowska
Elephant Man	http://en.wikipedia.org/wiki/Elephant_Man_(musician)
Elfriede Jelinek	http://en.wikipedia.org/wiki/Elfriede_Jelinek
Elfyn Llwyd	http://en.wikipedia.org/wiki/Elfyn_Llwyd
Elgin Baylor	http://en.wikipedia.org/wiki/Elgin_Baylor
Eli Jacobs	http://en.wikipedia.org/wiki/Eli_Jacobs
Eli Manning	http://en.wikipedia.org/wiki/Eli_Manning
Eli Wallach	http://en.wikipedia.org/wiki/Eli_Wallach
Eli Whitney	http://en.wikipedia.org/wiki/Eli_Whitney
Elia Kazan	http://en.wikipedia.org/wiki/Elia_Kazan
Elian Gonzalez	http://en.wikipedia.org/wiki/Elian_Gonzalez
Eliana Alexander	http://en.wikipedia.org/wiki/Eliana_Alexander
Elias Hicks	http://en.wikipedia.org/wiki/Elias_Hicks
Elias Howe	http://en.wikipedia.org/wiki/Elias_Howe
Elias James Corey	http://en.wikipedia.org/wiki/Elias_James_Corey
�lie Dot�	http://en.wikipedia.org/wiki/Elie_Dot%C3%A9
�lie Ducommun	http://en.wikipedia.org/wiki/%C9lie_Ducommun
�lie Faure	http://en.wikipedia.org/wiki/%C9lie_Faure
Elie Wiesel	http://en.wikipedia.org/wiki/Elie_Wiesel
Eliel Saarinen	http://en.wikipedia.org/wiki/Eliel_Saarinen
Elihu Benjamin Washburne	http://en.wikipedia.org/wiki/Elihu_Benjamin_Washburne
Elihu Burritt	http://en.wikipedia.org/wiki/Elihu_Burritt
Elihu Root	http://en.wikipedia.org/wiki/Elihu_Root
Elijah Cummings	http://en.wikipedia.org/wiki/Elijah_Cummings
Elijah Muhammad	http://en.wikipedia.org/wiki/Elijah_Muhammad
Elijah Wood	http://en.wikipedia.org/wiki/Elijah_Wood
Elinor Donahue	http://en.wikipedia.org/wiki/Elinor_Donahue
Elinor Wylie	http://en.wikipedia.org/wiki/Elinor_Wylie
Elio Vittorini	http://en.wikipedia.org/wiki/Elio_Vittorini
Eliot Engel	http://en.wikipedia.org/wiki/Eliot_Engel
Eliot Ness	http://en.wikipedia.org/wiki/Eliot_Ness
Eliot Spitzer	http://en.wikipedia.org/wiki/Eliot_Spitzer
Elisabeth Bumiller	http://en.wikipedia.org/wiki/Elisabeth_Bumiller
Elisabeth K�bler-Ross	http://en.wikipedia.org/wiki/Elisabeth_K%C3%BCbler-Ross
Elisabeth Moss	http://en.wikipedia.org/wiki/Elisabeth_Moss
Elisabeth Rohm	http://en.wikipedia.org/wiki/Elisabeth_Rohm
Elisabeth Shue	http://en.wikipedia.org/wiki/Elisabeth_Shue
Elisabeth Sladen	http://en.wikipedia.org/wiki/Elisabeth_Sladen
Elise Neal	http://en.wikipedia.org/wiki/Elise_Neal
Elisha Cuthbert	http://en.wikipedia.org/wiki/Elisha_Cuthbert
Eliza Dushku	http://en.wikipedia.org/wiki/Eliza_Dushku
Eliza Haywood	http://en.wikipedia.org/wiki/Eliza_Haywood
Elizabeth Alvarez	http://en.wikipedia.org/wiki/Elizabeth_Alvarez
Elizabeth Ashley	http://en.wikipedia.org/wiki/Elizabeth_Ashley
Elizabeth Báthory	http://en.wikipedia.org/wiki/Elizabeth_B%C3%A1thory
Elizabeth Barrett Browning	http://en.wikipedia.org/wiki/Elizabeth_Barrett_Browning
Elizabeth Berkley	http://en.wikipedia.org/wiki/Elizabeth_Berkley
Elizabeth Bishop	http://en.wikipedia.org/wiki/Elizabeth_Bishop
Elizabeth Bowen	http://en.wikipedia.org/wiki/Elizabeth_Bowen
Elizabeth Bowes-Lyon	http://en.wikipedia.org/wiki/Elizabeth_Bowes-Lyon
Elizabeth Burkley	http://en.wikipedia.org/wiki/Elizabeth_Berkley
Elizabeth Cady Stanton	http://en.wikipedia.org/wiki/Elizabeth_Cady_Stanton
Elizabeth Clare Prophet	http://en.wikipedia.org/wiki/Elizabeth_Clare_Prophet
Elizabeth Cleghorn Gaskell	http://en.wikipedia.org/wiki/Elizabeth_Cleghorn_Gaskell
Elizabeth Daily	http://en.wikipedia.org/wiki/Elizabeth_Daily
Elizabeth Dole	http://en.wikipedia.org/wiki/Elizabeth_Dole
Elizabeth Drew	http://en.wikipedia.org/wiki/Elizabeth_Drew
Elizabeth Fraser	http://en.wikipedia.org/wiki/Elizabeth_Fraser
Elizabeth Gracen	http://en.wikipedia.org/wiki/Elizabeth_Gracen
Elizabeth Hardwick	http://en.wikipedia.org/wiki/Elizabeth_Hardwick_(writer)
Elizabeth Hurley	http://en.wikipedia.org/wiki/Elizabeth_Hurley
Elizabeth II	http://en.wikipedia.org/wiki/Elizabeth_II
Elizabeth II	http://en.wikipedia.org/wiki/Elizabeth_II
Elizabeth II	http://en.wikipedia.org/wiki/Elizabeth_II
Elizabeth II	http://en.wikipedia.org/wiki/Elizabeth_II
Elizabeth II	http://en.wikipedia.org/wiki/Elizabeth_II
Elizabeth II	http://en.wikipedia.org/wiki/Elizabeth_II
Elizabeth II	http://en.wikipedia.org/wiki/Elizabeth_II
Elizabeth II	http://en.wikipedia.org/wiki/Elizabeth_II
Elizabeth II	http://en.wikipedia.org/wiki/Elizabeth_II
Elizabeth II	http://en.wikipedia.org/wiki/Elizabeth_II
Elizabeth II	http://en.wikipedia.org/wiki/Elizabeth_II
Elizabeth II	http://en.wikipedia.org/wiki/Elizabeth_II
Elizabeth II	http://en.wikipedia.org/wiki/Elizabeth_II
Elizabeth II	http://en.wikipedia.org/wiki/Elizabeth_II
Elizabeth II	http://en.wikipedia.org/wiki/Elizabeth_II
Elizabeth II	http://en.wikipedia.org/wiki/Elizabeth_II
Elizabeth II	http://en.wikipedia.org/wiki/Elizabeth_II
Elizabeth II	http://en.wikipedia.org/wiki/Elizabeth_II
Elizabeth II	http://en.wikipedia.org/wiki/Elizabeth_II
Elizabeth Jennings	http://en.wikipedia.org/wiki/Elizabeth_Jennings
Elizabeth Jolley	http://en.wikipedia.org/wiki/Elizabeth_Jolley
Elizabeth Kendall	http://en.wikipedia.org/wiki/Elizabeth_Kendall
Elizabeth Madox Roberts	http://en.wikipedia.org/wiki/Elizabeth_Madox_Roberts
Elizabeth McGovern	http://en.wikipedia.org/wiki/Elizabeth_McGovern
Elizabeth Mitchell	http://en.wikipedia.org/wiki/Elizabeth_Mitchell
Elizabeth Montagu	http://en.wikipedia.org/wiki/Elizabeth_Montagu
Elizabeth Montgomery	http://en.wikipedia.org/wiki/Elizabeth_Montgomery
Elizabeth Moon	http://en.wikipedia.org/wiki/Elizabeth_Moon
Elizabeth Pe�a	http://en.wikipedia.org/wiki/Elizabeth_Pe%C3%B1a
Elizabeth Perkins	http://en.wikipedia.org/wiki/Elizabeth_Perkins
Elizabeth Sanderson Haldane	http://en.wikipedia.org/wiki/Elizabeth_Sanderson_Haldane
Elizabeth Smart	http://en.wikipedia.org/wiki/Elizabeth_Smart_%28activist%29
Elizabeth Stuart Phelps Ward	http://en.wikipedia.org/wiki/Elizabeth_Stuart_Phelps_Ward
Elizabeth Taylor	http://en.wikipedia.org/wiki/Elizabeth_Taylor
Elizabeth Truss	http://en.wikipedia.org/wiki/Elizabeth_Truss
Elizabeth Vargas	http://en.wikipedia.org/wiki/Elizabeth_Vargas
Elizabeth Warren	http://en.wikipedia.org/wiki/Elizabeth_Warren
Elizebeth Friedman	http://en.wikipedia.org/wiki/Elizebeth_Friedman
Elke Sommer	http://en.wikipedia.org/wiki/Elke_Sommer
Ella Fitzgerald	http://en.wikipedia.org/wiki/Ella_Fitzgerald
Ella T. Grasso	http://en.wikipedia.org/wiki/Ella_T._Grasso
Ella Wheeler Wilcox	http://en.wikipedia.org/wiki/Ella_Wheeler_Wilcox
Elle Fanning	http://en.wikipedia.org/wiki/Elle_Fanning
Elle Macpherson	http://en.wikipedia.org/wiki/Elle_Macpherson
Ellen Albertini Dow	http://en.wikipedia.org/wiki/Ellen_Albertini_Dow
Ellen Barkin	http://en.wikipedia.org/wiki/Ellen_Barkin
Ellen Burstyn	http://en.wikipedia.org/wiki/Ellen_Burstyn
Ellen Corby	http://en.wikipedia.org/wiki/Ellen_Corby
Ellen DeGeneres	http://en.wikipedia.org/wiki/Ellen_DeGeneres
Ellen Drew	http://en.wikipedia.org/wiki/Ellen_Drew
Ellen Feiss	http://en.wikipedia.org/wiki/Ellen_Feiss
Ellen G. White	http://en.wikipedia.org/wiki/Ellen_G._White
Ellen Gilchrist	http://en.wikipedia.org/wiki/Ellen_Gilchrist
Ellen Glasgow	http://en.wikipedia.org/wiki/Ellen_Glasgow
Ellen Goodman	http://en.wikipedia.org/wiki/Ellen_Goodman
Ellen Johnson-Sirleaf	http://en.wikipedia.org/wiki/Ellen_Johnson-Sirleaf
Ellen Malcolm	http://en.wikipedia.org/wiki/Ellen_Malcolm
Ellen Muth	http://en.wikipedia.org/wiki/Ellen_Muth
Ellen Pompeo	http://en.wikipedia.org/wiki/Ellen_Pompeo
Ellen Tauscher	http://en.wikipedia.org/wiki/Ellen_Tauscher
Elliot Richardson	http://en.wikipedia.org/wiki/Elliot_Richardson
Elliot Sharp	http://en.wikipedia.org/wiki/Elliott_Sharp
Elliott Abrams	http://en.wikipedia.org/wiki/Elliott_Abrams
Elliott Baker	http://en.wikipedia.org/wiki/Elliott_Baker
Elliott Carter	http://en.wikipedia.org/wiki/Elliott_Carter
Elliott Gould	http://en.wikipedia.org/wiki/Elliott_Gould
Elliott Murphy	http://en.wikipedia.org/wiki/Elliott_Murphy
Elliott Smith	http://en.wikipedia.org/wiki/Elliott_Smith
Elmer Bernstein	http://en.wikipedia.org/wiki/Elmer_Bernstein
Elmer Rice	http://en.wikipedia.org/wiki/Elmer_Rice
Elmer Wayne Henley	http://en.wikipedia.org/wiki/Elmer_Wayne_Henley
Elmo Roper	http://en.wikipedia.org/wiki/Elmo_Roper
Elmore Leonard	http://en.wikipedia.org/wiki/Elmore_Leonard
Elpidio Quirino	http://en.wikipedia.org/wiki/Elpidio_Quirino
Elroy "Crazy Legs" Hirsch	http://en.wikipedia.org/wiki/Elroy_%22Crazy_Legs%22_Hirsch
Elsa Lanchester	http://en.wikipedia.org/wiki/Elsa_Lanchester
Elsa Martinelli	http://en.wikipedia.org/wiki/Elsa_Martinelli
Elton Gallegly	http://en.wikipedia.org/wiki/Elton_Gallegly
Elton John	http://en.wikipedia.org/wiki/Elton_John
Elvin Bishop	http://en.wikipedia.org/wiki/Elvin_Bishop
Elvin Jones	http://en.wikipedia.org/wiki/Elvin_Jones
Elvis Costello	http://en.wikipedia.org/wiki/Elvis_Costello
Elvis Mitchell	http://en.wikipedia.org/wiki/Elvis_Mitchell
Elvis Presley	http://en.wikipedia.org/wiki/Elvis_Presley
Elwood Hillis	http://en.wikipedia.org/wiki/Elwood_Hillis
Ely Ould Mohamed Vall	http://en.wikipedia.org/wiki/Ely_Ould_Mohamed_Vall
Emanuel Bronner	http://en.wikipedia.org/wiki/Emanuel_Bronner
Emanuel Cleaver	http://en.wikipedia.org/wiki/Emanuel_Cleaver
Emanuel Swedenborg	http://en.wikipedia.org/wiki/Emanuel_Swedenborg
Emelian Pugachev	http://en.wikipedia.org/wiki/Emelian_Pugachev
Emeric Pressburger	http://en.wikipedia.org/wiki/Emeric_Pressburger
Emeril Lagasse	http://en.wikipedia.org/wiki/Emeril_Lagasse
Emerson Fittipaldi	http://en.wikipedia.org/wiki/Emerson_Fittipaldi
Emil Boc	http://en.wikipedia.org/wiki/Emil_Boc
Emil Fischer	http://en.wikipedia.org/wiki/Hermann_Emil_Fischer
Emil Jannings	http://en.wikipedia.org/wiki/Emil_Jannings
Emil Ludwig	http://en.wikipedia.org/wiki/Emil_Ludwig
Emil von Behring	http://en.wikipedia.org/wiki/Emil_von_Behring
�mile Durkheim	http://en.wikipedia.org/wiki/%C9mile_Durkheim
Emile Hirsch	http://en.wikipedia.org/wiki/Emile_Hirsch
Emile Lahoud	http://en.wikipedia.org/wiki/Emile_Lahoud
�mile Zola	http://en.wikipedia.org/wiki/%C9mile_Zola
Emiliano Zapata	http://en.wikipedia.org/wiki/Emiliano_Zapata
Emilie de Ravin	http://en.wikipedia.org/wiki/Emilie_de_Ravin
Emilie Dionne	http://en.wikipedia.org/wiki/Dionne_quintuplets
Emilinha Borba	http://en.wikipedia.org/wiki/Emilinha_Borba
Emilio Aguinaldo	http://en.wikipedia.org/wiki/Emilio_Aguinaldo
Emilio Estevez	http://en.wikipedia.org/wiki/Emilio_Estevez
Emilio G. Segr�	http://en.wikipedia.org/wiki/Emilio_Segr%C3%A8
Emilio Garza	http://en.wikipedia.org/wiki/Emilio_Garza
Emily Anne Eliza Shirreff	http://en.wikipedia.org/wiki/Emily_Anne_Eliza_Shirreff
Emily Bront�	http://en.wikipedia.org/wiki/Emily_Bront%C3%AB
Emily Browning	http://en.wikipedia.org/wiki/Emily_Browning
Emily Carter	http://en.wikipedia.org/wiki/Emily_Carter
Emily de Jongh-Elhage	http://en.wikipedia.org/wiki/Emily_de_Jongh-Elhage
Emily Dickinson	http://en.wikipedia.org/wiki/Emily_Dickinson
Emily Greene Balch	http://en.wikipedia.org/wiki/Emily_Greene_Balch
Emily Lloyd	http://en.wikipedia.org/wiki/Emily_Lloyd
Emily Mortimer	http://en.wikipedia.org/wiki/Emily_Mortimer
Emily Post	http://en.wikipedia.org/wiki/Emily_Post
Emily Procter	http://en.wikipedia.org/wiki/Emily_Procter
Emily Saliers	http://en.wikipedia.org/wiki/Emily_Saliers
Emily Thornberry	http://en.wikipedia.org/wiki/Emily_Thornberry
Emily VanCamp	http://en.wikipedia.org/wiki/Emily_VanCamp
Emily Watson	http://en.wikipedia.org/wiki/Emily_Watson
Emin Pasha	http://en.wikipedia.org/wiki/Emin_Pasha
Emir Kusturica	http://en.wikipedia.org/wiki/Emir_Kusturica
Emma Anderson	http://en.wikipedia.org/wiki/Emma_Anderson
Emma Bunton	http://en.wikipedia.org/wiki/Emma_Bunton
Emma Goldman	http://en.wikipedia.org/wiki/Emma_Goldman
Emma Hamilton	http://en.wikipedia.org/wiki/Emma_Hamilton
Emma Lazarus	http://en.wikipedia.org/wiki/Emma_Lazarus
Emma Reynolds	http://en.wikipedia.org/wiki/Emma_Reynolds
Emma Roberts	http://en.wikipedia.org/wiki/Emma_Roberts
Emma Samms	http://en.wikipedia.org/wiki/Emma_Samms
Emma Thompson	http://en.wikipedia.org/wiki/Emma_Thompson
Emma Watson	http://en.wikipedia.org/wiki/Emma_Watson
Emmanuel Goldstein	http://en.wikipedia.org/wiki/Emmanuel_Goldstein
Emmanuel Levinas	http://en.wikipedia.org/wiki/Emmanuel_Levinas
Emmanuel Lewis	http://en.wikipedia.org/wiki/Emmanuel_Lewis
Emmanuel Nadingar	http://en.wikipedia.org/wiki/Emmanuel_Nadingar
Emmanuel Philibert	http://en.wikipedia.org/wiki/Emmanuel_Philibert
Emmanuelle B�art	http://en.wikipedia.org/wiki/Emmanuelle_B%C3%A9art
Emmeline Pankhurst	http://en.wikipedia.org/wiki/Emmeline_Pankhurst
Emmett Till	http://en.wikipedia.org/wiki/Emmett_Till
Emmitt Smith	http://en.wikipedia.org/wiki/Emmitt_Smith
Emmy Rossum	http://en.wikipedia.org/wiki/Emmy_Rossum
Emmylou Harris	http://en.wikipedia.org/wiki/Emmylou_Harris
Emo Philips	http://en.wikipedia.org/wiki/Emo_Philips
Emomalii Rahmon	http://en.wikipedia.org/wiki/Emomalii_Rahmon
Emperor Akihito	http://en.wikipedia.org/wiki/Emperor_Akihito
Emperor Bokassa I	http://en.wikipedia.org/wiki/Jean-B%C3%A9del_Bokassa
Emperor Hirohito	http://en.wikipedia.org/wiki/Emperor_Hirohito
Emperor Norton	http://en.wikipedia.org/wiki/Emperor_Norton
Empress Michiko	http://en.wikipedia.org/wiki/Empress_Michiko
Engelbert Humperdinck	http://en.wikipedia.org/wiki/Engelbert_Humperdinck
Eni Faleomavaega	http://en.wikipedia.org/wiki/Eni_Faleomavaega
Enid Bagnold	http://en.wikipedia.org/wiki/Enid_Bagnold
Ennio Morricone	http://en.wikipedia.org/wiki/Ennio_Morricone
Enoch Powell	http://en.wikipedia.org/wiki/Enoch_Powell
Enos T. Throop	http://en.wikipedia.org/wiki/Enos_T._Throop
Enrico Caruso	http://en.wikipedia.org/wiki/Enrico_Caruso
Enrico Fermi	http://en.wikipedia.org/wiki/Enrico_Fermi
Enrique Bola�os	http://en.wikipedia.org/wiki/Enrique_Bola%C3%B1os
Enrique Granados	http://en.wikipedia.org/wiki/Enrique_Granados
Enrique Iglesias	http://en.wikipedia.org/wiki/Enrique_Iglesias
Enver Hoxha	http://en.wikipedia.org/wiki/Enver_Hoxha
Enver Pasha	http://en.wikipedia.org/wiki/Enver_Pasha
Enzo Ferrari	http://en.wikipedia.org/wiki/Enzo_Ferrari
Epeli Nailatikau	http://en.wikipedia.org/wiki/Epeli_Nailatikau
Ephraim Chambers	http://en.wikipedia.org/wiki/Ephraim_Chambers
Ephraim Inoni	http://en.wikipedia.org/wiki/Ephraim_Inoni
Erasmus Alberus	http://en.wikipedia.org/wiki/Erasmus_Alberus
Erasmus Darwin	http://en.wikipedia.org/wiki/Erasmus_Darwin
Eric A. Cornell	http://en.wikipedia.org/wiki/Eric_A._Cornell
Eric Alterman	http://en.wikipedia.org/wiki/Eric_Alterman
Eric Ambler	http://en.wikipedia.org/wiki/Eric_Ambler
Eric Andersen	http://en.wikipedia.org/wiki/Eric_Andersen
Eric Avery	http://en.wikipedia.org/wiki/Eric_Avery
Eric Balfour	http://en.wikipedia.org/wiki/Eric_Balfour
Eric Bana	http://en.wikipedia.org/wiki/Eric_Bana
Eric Ben�t	http://en.wikipedia.org/wiki/Eric_Ben%C3%A9t
Eric Bentley	http://en.wikipedia.org/wiki/Eric_Bentley
Eric Bogosian	http://en.wikipedia.org/wiki/Eric_Bogosian
Eric Braeden	http://en.wikipedia.org/wiki/Eric_Braeden
Eric Burdon	http://en.wikipedia.org/wiki/Eric_Burdon
Eric Burns	http://en.wikipedia.org/wiki/Eric_Burns
Eric Cantona	http://en.wikipedia.org/wiki/Eric_Cantona
Eric Cantor	http://en.wikipedia.org/wiki/Eric_Cantor
Eric Carr	http://en.wikipedia.org/wiki/Eric_Carr
Eric Christian Olsen	http://en.wikipedia.org/wiki/Eric_Christian_Olsen
Eric Clapton	http://en.wikipedia.org/wiki/Eric_Clapton
Eric Close	http://en.wikipedia.org/wiki/Eric_Close
Eric Dolphy	http://en.wikipedia.org/wiki/Eric_Dolphy
Eric Erlandson	http://en.wikipedia.org/wiki/Eric_Erlandson
Eric Gill	http://en.wikipedia.org/wiki/Eric_Gill
Eric Harris	http://en.wikipedia.org/wiki/Eric_David_Harris
Eric Heiden	http://en.wikipedia.org/wiki/Eric_Heiden
Eric Hoffer	http://en.wikipedia.org/wiki/Eric_Hoffer
Eric Holder	http://en.wikipedia.org/wiki/Eric_Holder
Eric Idle	http://en.wikipedia.org/wiki/Eric_Idle
Eric Idle	http://en.wikipedia.org/wiki/Eric_Idle
Eric Illsley	http://en.wikipedia.org/wiki/Eric_Illsley
Eric Johnson	http://en.wikipedia.org/wiki/Eric_Johnson_(actor)
Eric Johnson	http://en.wikipedia.org/wiki/Eric_Johnson
Eric Joyce	http://en.wikipedia.org/wiki/Eric_Joyce
Eric Lichtblau	http://en.wikipedia.org/wiki/Eric_Lichtblau
Eric Lindros	http://en.wikipedia.org/wiki/Eric_Lindros
Eric Lloyd	http://en.wikipedia.org/wiki/Eric_Lloyd
Eric Lutes	http://en.wikipedia.org/wiki/Eric_Lutes
Eric Mabius	http://en.wikipedia.org/wiki/Eric_Mabius
Eric McCormack	http://en.wikipedia.org/wiki/Eric_McCormack
Eric Morecambe	http://en.wikipedia.org/wiki/Eric_Morecambe
Eric Ollerenshaw	http://en.wikipedia.org/wiki/Eric_Ollerenshaw
Eric Pickles	http://en.wikipedia.org/wiki/Eric_Pickles
Eric Roberts	http://en.wikipedia.org/wiki/Eric_Roberts
�ric Rohmer	http://en.wikipedia.org/wiki/%C9ric_Rohmer
Eric Rudolph	http://en.wikipedia.org/wiki/Eric_Rudolph
Eric S. Raymond	http://en.wikipedia.org/wiki/Eric_S._Raymond
Eric Schmidt	http://en.wikipedia.org/wiki/Eric_Schmidt
Eric Sevareid	http://en.wikipedia.org/wiki/Eric_Sevareid
Eric Shinseki	http://en.wikipedia.org/wiki/Eric_Shinseki
Eric Stefani	http://en.wikipedia.org/wiki/Eric_Stefani
Eric Stewart	http://en.wikipedia.org/wiki/Eric_Stewart
Eric Stoltz	http://en.wikipedia.org/wiki/Eric_Stoltz
Eric Szmanda	http://en.wikipedia.org/wiki/Eric_Szmanda
Eric Walrond	http://en.wikipedia.org/wiki/Eric_Walrond
Eric Woolfson	http://en.wikipedia.org/wiki/Eric_Woolfson
Erica Durance	http://en.wikipedia.org/wiki/Erica_Durance
Erica Gavin	http://en.wikipedia.org/wiki/Erica_Gavin
Erica Jong	http://en.wikipedia.org/wiki/Erica_Jong
Erich Fromm	http://en.wikipedia.org/wiki/Erich_Fromm
Erich Honecker	http://en.wikipedia.org/wiki/Erich_Honecker
Erich Maria Remarque	http://en.wikipedia.org/wiki/Erich_Maria_Remarque
Erich Raeder	http://en.wikipedia.org/wiki/Erich_Raeder
Erich Topp	http://en.wikipedia.org/wiki/Erich_Topp
Erich von D�niken	http://en.wikipedia.org/wiki/Erich_von_D%C3%A4niken
Erich von Manstein	http://en.wikipedia.org/wiki/Erich_von_Manstein
Erich von Stroheim	http://en.wikipedia.org/wiki/Erich_von_Stroheim
Erik Aaes	http://en.wikipedia.org/wiki/Erik_Aaes
Erik Aud�	http://en.wikipedia.org/wiki/Erik_Aud%C3%A9
Erik Erikson	http://en.wikipedia.org/wiki/Erik_Erikson
Erik Estrada	http://en.wikipedia.org/wiki/Erik_Estrada
Erik Fleming	http://en.wikipedia.org/wiki/Erik_Fleming_(director)
Erik Menendez	http://en.wikipedia.org/wiki/Erik_Menendez
Erik Paulsen	http://en.wikipedia.org/wiki/Erik_Paulsen
Erik Prince	http://en.wikipedia.org/wiki/Erik_Prince
Erik Satie	http://en.wikipedia.org/wiki/Erik_Satie
Erik von Detten	http://en.wikipedia.org/wiki/Erik_von_Detten
Erik von Kuehnelt-Leddihn	http://en.wikipedia.org/wiki/Erik_von_Kuehnelt-Leddihn
Erik XIV	http://en.wikipedia.org/wiki/Erik_XIV
Erika Alexander	http://en.wikipedia.org/wiki/Erika_Alexander
Erika Christensen	http://en.wikipedia.org/wiki/Erika_Christensen
Erika Eleniak	http://en.wikipedia.org/wiki/Erika_Eleniak
Erika Mann	http://en.wikipedia.org/wiki/Erika_Mann
Erika Slezak	http://en.wikipedia.org/wiki/Erika_Slezak
Erin Brockovich	http://en.wikipedia.org/wiki/Erin_Brockovich
Erin Daniels	http://en.wikipedia.org/wiki/Erin_Daniels
Erin Gray	http://en.wikipedia.org/wiki/Erin_Gray
Erin Moran	http://en.wikipedia.org/wiki/Erin_Moran
Eriq La Salle	http://en.wikipedia.org/wiki/Eriq_La_Salle
Erle Stanley Gardner	http://en.wikipedia.org/wiki/Erle_Stanley_Gardner
Erma Bombeck	http://en.wikipedia.org/wiki/Erma_Bombeck
Ermanno Olmi	http://en.wikipedia.org/wiki/Ermanno_Olmi
Ernest Bai Koroma	http://en.wikipedia.org/wiki/Ernest_Bai_Koroma
Ernest Bloch	http://en.wikipedia.org/wiki/Ernest_Bloch
Ernest Borgnine	http://en.wikipedia.org/wiki/Ernest_Borgnine
Ernest Buckler	http://en.wikipedia.org/wiki/Ernest_Buckler
Ernest Burgess	http://en.wikipedia.org/wiki/Ernest_Burgess
Ernest Dowson	http://en.wikipedia.org/wiki/Ernest_Dowson
Ernest F. Hollings	http://en.wikipedia.org/wiki/Ernest_F._Hollings
Ernest Gallo	http://en.wikipedia.org/wiki/Gallo_family
Ernest Gruening	http://en.wikipedia.org/wiki/Ernest_Gruening
Ernest Hemingway	http://en.wikipedia.org/wiki/Ernest_Hemingway
Ernest Istook	http://en.wikipedia.org/wiki/Ernest_Istook
Ernest Lawrence	http://en.wikipedia.org/wiki/Ernest_Lawrence
Ernest Poole	http://en.wikipedia.org/wiki/Ernest_Poole
Ernest Rutherford	http://en.wikipedia.org/wiki/Ernest_Rutherford
Ernest T. S. Walton	http://en.wikipedia.org/wiki/Ernest_Walton
Ernest Thesiger	http://en.wikipedia.org/wiki/Ernest_Thesiger
Ernest Tubb	http://en.wikipedia.org/wiki/Ernest_Tubb
Ernest van den Haag	http://en.wikipedia.org/wiki/Ernest_van_den_Haag
Ernesto Cardenal	http://en.wikipedia.org/wiki/Ernesto_Cardenal
Ernesto Sábato	http://en.wikipedia.org/wiki/Ernesto_S%C3%A1bato
Ernesto Teodoro Moneta	http://en.wikipedia.org/wiki/Ernesto_Teodoro_Moneta
Ernesto Zedillo	http://en.wikipedia.org/wiki/Ernesto_Zedillo
Ernie Banks	http://en.wikipedia.org/wiki/Ernie_Banks
Ernie Fletcher	http://en.wikipedia.org/wiki/Ernie_Fletcher
Ernie Fletcher	http://en.wikipedia.org/wiki/Ernie_Fletcher
Ernie Harwell	http://en.wikipedia.org/wiki/Ernie_Harwell
Ernie Hudson	http://en.wikipedia.org/wiki/Ernie_Hudson
Ernie Kovacs	http://en.wikipedia.org/wiki/Ernie_Kovacs
Ernie Pyle	http://en.wikipedia.org/wiki/Ernie_Pyle
Ernie Wise	http://en.wikipedia.org/wiki/Ernie_Wise
Erno Rubik	http://en.wikipedia.org/wiki/Erno_Rubik
Ernst Engel	http://en.wikipedia.org/wiki/Ernst_Engel
Ernst Haeckel	http://en.wikipedia.org/wiki/Ernst_Haeckel
Ernst Kaltenbrunner	http://en.wikipedia.org/wiki/Ernst_Kaltenbrunner
Ernst Lubitsch	http://en.wikipedia.org/wiki/Ernst_Lubitsch
Ernst Mach	http://en.wikipedia.org/wiki/Ernst_Mach
Ernst Mayr	http://en.wikipedia.org/wiki/Ernst_Mayr
Ernst Otto Fischer	http://en.wikipedia.org/wiki/Ernst_Otto_Fischer
Ernst Roehm	http://en.wikipedia.org/wiki/Ernst_Roehm
Ernst Ruska	http://en.wikipedia.org/wiki/Ernst_Ruska
Ernst Winar	http://en.wikipedia.org/wiki/Ernst_Winar
Ernst Zundel	http://en.wikipedia.org/wiki/Ernst_Zundel
Errol Braithwaite	http://en.wikipedia.org/wiki/Errol_Braithwaite
Errol Flynn	http://en.wikipedia.org/wiki/Errol_Flynn
Errol Morris	http://en.wikipedia.org/wiki/Errol_Morris
Erskine Bowles	http://en.wikipedia.org/wiki/Erskine_Bowles
Erskine Caldwell	http://en.wikipedia.org/wiki/Erskine_Caldwell
Ervin Drake	http://en.wikipedia.org/wiki/Ervin_Drake
Erving Goffman	http://en.wikipedia.org/wiki/Erving_Goffman
Erwin Rommel	http://en.wikipedia.org/wiki/Erwin_Rommel
Erwin Schr�dinger	http://en.wikipedia.org/wiki/Erwin_Schr%C3%B6dinger
Erwin von Witzleben	http://en.wikipedia.org/wiki/Erwin_von_Witzleben
Erykah Badu	http://en.wikipedia.org/wiki/Erykah_Badu
Esai Morales	http://en.wikipedia.org/wiki/Esai_Morales
Esaias Tegn�r	http://en.wikipedia.org/wiki/Esaias_Tegn%C3%A9r
Esa-Pekka Salonen	http://en.wikipedia.org/wiki/Esa-Pekka_Salonen
Essie Mae Washington-Williams	http://en.wikipedia.org/wiki/Essie_Mae_Washington-Williams
Esteban E. Torres	http://en.wikipedia.org/wiki/Esteban_E._Torres
Est�e Lauder	http://en.wikipedia.org/wiki/Est%C3%A9e_Lauder_%28person%29
Estella Warren	http://en.wikipedia.org/wiki/Estella_Warren
Estelle Getty	http://en.wikipedia.org/wiki/Estelle_Getty
Estelle Parsons	http://en.wikipedia.org/wiki/Estelle_Parsons
Estelle Winwood	http://en.wikipedia.org/wiki/Estelle_Winwood
Estes Kefauver	http://en.wikipedia.org/wiki/Estes_Kefauver
Esther Dyson	http://en.wikipedia.org/wiki/Esther_Dyson
Esther McVey	http://en.wikipedia.org/wiki/Esther_McVey
Esther Rolle	http://en.wikipedia.org/wiki/Esther_Rolle
Esther Williams	http://en.wikipedia.org/wiki/Esther_Williams
Ethan Allen	http://en.wikipedia.org/wiki/Ethan_Allen
Ethan Coen	http://en.wikipedia.org/wiki/Ethan_Coen
Ethan Embry	http://en.wikipedia.org/wiki/Ethan_Embry
Ethan Hawke	http://en.wikipedia.org/wiki/Ethan_Hawke
Ethan Suplee	http://en.wikipedia.org/wiki/Ethan_Suplee
Ethel Barrymore	http://en.wikipedia.org/wiki/Ethel_Barrymore
Ethel Kennedy	http://en.wikipedia.org/wiki/Ethel_Kennedy
Ethel Mannin	http://en.wikipedia.org/wiki/Ethel_Mannin
Ethel Merman	http://en.wikipedia.org/wiki/Ethel_Merman
Ethel Rosenberg	http://en.wikipedia.org/wiki/Ethel_Rosenberg
Ethel Waters	http://en.wikipedia.org/wiki/Ethel_Waters
Etheridge Knight	http://en.wikipedia.org/wiki/Etheridge_Knight
�tienne Louis Malus	http://en.wikipedia.org/wiki/%C9tienne_Louis_Malus
�tienne Pasquier	http://en.wikipedia.org/wiki/%C9tienne_Pasquier
Etienne Ys	http://en.wikipedia.org/wiki/Etienne_Ys
�tienne-Denis Pasquier	http://en.wikipedia.org/wiki/%C9tienne-Denis_Pasquier
Etta James	http://en.wikipedia.org/wiki/Etta_James
Eubie Blake	http://en.wikipedia.org/wiki/Eubie_Blake
Eudora Welty	http://en.wikipedia.org/wiki/Eudora_Welty
Eudoxus of Cnidus	http://en.wikipedia.org/wiki/Eudoxus_of_Cnidus
Eugen Bleuler	http://en.wikipedia.org/wiki/Eugen_Bleuler
Eugen Weber	http://en.wikipedia.org/wiki/Eugen_Weber
Eugene A. Chappie	http://en.wikipedia.org/wiki/Eugene_A._Chappie
Eugene Allen	http://en.wikipedia.org/wiki/Robert_Eugene_Allen
Eugene Asa Carr	http://en.wikipedia.org/wiki/Eugene_Asa_Carr
Eugene Chadbourne	http://en.wikipedia.org/wiki/Eugene_Chadbourne
Eug�ne Delacroix	http://en.wikipedia.org/wiki/Eug%C3%A8ne_Delacroix
Eugene Field	http://en.wikipedia.org/wiki/Eugene_Field
Eug�ne Ionesco	http://en.wikipedia.org/wiki/Eug%C3%A8ne_Ionesco
Eugene Jolas	http://en.wikipedia.org/wiki/Eugene_Jolas
Eugene Levy	http://en.wikipedia.org/wiki/Eugene_Levy
Eugene Lyons	http://en.wikipedia.org/wiki/Eugene_Lyons
Eugene McCarthy	http://en.wikipedia.org/wiki/Eugene_McCarthy
Eugene Meyer	http://en.wikipedia.org/wiki/Eugene_Meyer
Eugene O. Sykes	http://en.wikipedia.org/wiki/Eugene_O._Sykes
Eugene O'Neill	http://en.wikipedia.org/wiki/Eugene_O%27Neill
Eugene R. McGrath	http://en.wikipedia.org/wiki/Eugene_R._McGrath
Eug�ne Sue	http://en.wikipedia.org/wiki/Eug%C3%A8ne_Sue
Eugene V. Debs	http://en.wikipedia.org/wiki/Eugene_V._Debs
Eugene Wigner	http://en.wikipedia.org/wiki/Eugene_Wigner
Eugenie Anderson	http://en.wikipedia.org/wiki/Eugenie_Anderson
Eugenio Montale	http://en.wikipedia.org/wiki/Eugenio_Montale
Eunice Kennedy Shriver	http://en.wikipedia.org/wiki/Eunice_Kennedy_Shriver
Eusebio Ferreira da Silva	http://en.wikipedia.org/wiki/Eus%C3%A9bio
Eustace John	http://en.wikipedia.org/wiki/Eustace_John
Eustache Deschamps	http://en.wikipedia.org/wiki/Eustache_Deschamps
Eva Amurri	http://en.wikipedia.org/wiki/Eva_Amurri
Eva Braun	http://en.wikipedia.org/wiki/Eva_Braun
Eva Gabor	http://en.wikipedia.org/wiki/Eva_Gabor
Eva Green	http://en.wikipedia.org/wiki/Eva_Green
Eva Herzigova	http://en.wikipedia.org/wiki/Eva_Herzigova
Eva LaRue	http://en.wikipedia.org/wiki/Eva_LaRue
Eva Longoria	http://en.wikipedia.org/wiki/Eva_Longoria
Eva Marie Saint	http://en.wikipedia.org/wiki/Eva_Marie_Saint
Eva Mendes	http://en.wikipedia.org/wiki/Eva_Mendes
Eva Tamargo Lemus	http://en.wikipedia.org/wiki/Eva_Tamargo
Evan Bayh	http://en.wikipedia.org/wiki/Evan_Bayh
Evan Dando	http://en.wikipedia.org/wiki/Evan_Dando
Evan Farmer	http://en.wikipedia.org/wiki/Evan_Farmer
Evan Handler	http://en.wikipedia.org/wiki/Evan_Handler
Evan Hunter	http://en.wikipedia.org/wiki/Evan_Hunter
Evan Lurie	http://en.wikipedia.org/wiki/Evan_Lurie_%28composer%29
Evan Mecham	http://en.wikipedia.org/wiki/Evan_Mecham
Evan Parker	http://en.wikipedia.org/wiki/Evan_Parker
Evan Rachel Wood	http://en.wikipedia.org/wiki/Evan_Rachel_Wood
Evander Holyfield	http://en.wikipedia.org/wiki/Evander_Holyfield
Evangeline Lilly	http://en.wikipedia.org/wiki/Evangeline_Lilly
Evangelista Torricelli	http://en.wikipedia.org/wiki/Evangelista_Torricelli
Eve Arden	http://en.wikipedia.org/wiki/Eve_Arden
Eve Plumb	http://en.wikipedia.org/wiki/Eve_Plumb
Evel Knievel	http://en.wikipedia.org/wiki/Evel_Knievel
Evelyn Ankers	http://en.wikipedia.org/wiki/Evelyn_Ankers
Evelyn Brent	http://en.wikipedia.org/wiki/Evelyn_Brent
Evelyn De Morgan	http://en.wikipedia.org/wiki/Evelyn_De_Morgan
Evelyn Glennie	http://en.wikipedia.org/wiki/Evelyn_Glennie
Evelyn Waugh	http://en.wikipedia.org/wiki/Evelyn_Waugh
Everett Dirksen	http://en.wikipedia.org/wiki/Everett_Dirksen
Everett McGill	http://en.wikipedia.org/wiki/Everett_McGill
Everett Sanders	http://en.wikipedia.org/wiki/Everett_Sanders
Everett Sloane	http://en.wikipedia.org/wiki/Everett_Sloane
Evgeny Baratynsky	http://en.wikipedia.org/wiki/Evgeny_Baratynsky
Evita Peron	http://en.wikipedia.org/wiki/Evita_Peron
Evo Morales	http://en.wikipedia.org/wiki/Evo_Morales
Evonne Goolagong	http://en.wikipedia.org/wiki/Evonne_Goolagong
Ewan McGregor	http://en.wikipedia.org/wiki/Ewan_McGregor
Exene Cervenka	http://en.wikipedia.org/wiki/Exene_Cervenka
Eydie Gorme	http://en.wikipedia.org/wiki/Eydie_Gorme
Ezer Weizman	http://en.wikipedia.org/wiki/Ezer_Weizman
Ezra Pound	http://en.wikipedia.org/wiki/Ezra_Pound
F. A. Hayek	http://en.wikipedia.org/wiki/F._A._Hayek
F. Donald Nixon	http://en.wikipedia.org/wiki/F._Donald_Nixon
F. H. Bradley	http://en.wikipedia.org/wiki/F._H._Bradley
F. James Sensenbrenner, Jr.	http://en.wikipedia.org/wiki/F._James_Sensenbrenner%2C_Jr.
F. Lee Bailey	http://en.wikipedia.org/wiki/F._Lee_Bailey
F. Marion Crawford	http://en.wikipedia.org/wiki/F._Marion_Crawford
F. Murray Abraham	http://en.wikipedia.org/wiki/F._Murray_Abraham
F. O. Matthiessen	http://en.wikipedia.org/wiki/F._O._Matthiessen
F. Scott Fitzgerald	http://en.wikipedia.org/wiki/F._Scott_Fitzgerald
F. Sherwood Rowland	http://en.wikipedia.org/wiki/F._Sherwood_Rowland
F. W. de Klerk	http://en.wikipedia.org/wiki/F._W._de_Klerk
Fabian Hamilton	http://en.wikipedia.org/wiki/Fabian_Hamilton
Fabio Capello	http://en.wikipedia.org/wiki/Fabio_Capello
Fabio Lanzoni	http://en.wikipedia.org/wiki/Fabio_Lanzoni
Fabrice Morvan	http://en.wikipedia.org/wiki/Fabrice_Morvan
Fabrizio Moretti	http://en.wikipedia.org/wiki/Fabrizio_Moretti
Fairuza Balk	http://en.wikipedia.org/wiki/Fairuza_Balk
Faisal I	http://en.wikipedia.org/wiki/Faisal_I
Faith Addis	http://en.wikipedia.org/wiki/Down_to_Earth_%28UK_TV_series%29
Faith Domergue	http://en.wikipedia.org/wiki/Faith_Domergue
Faith Evans	http://en.wikipedia.org/wiki/Faith_Evans
Faith Ford	http://en.wikipedia.org/wiki/Faith_Ford
Faith Hill	http://en.wikipedia.org/wiki/Faith_Hill
Famke Janssen	http://en.wikipedia.org/wiki/Famke_Janssen
Fannie Flagg	http://en.wikipedia.org/wiki/Fannie_Flagg
Fanny Ardant	http://en.wikipedia.org/wiki/Fanny_Ardant
Fanny Burney	http://en.wikipedia.org/wiki/Fanny_Burney
Fantasia Barrino	http://en.wikipedia.org/wiki/Fantasia_Barrino
Fareed Zakaria	http://en.wikipedia.org/wiki/Fareed_Zakaria
Farley Granger	http://en.wikipedia.org/wiki/Farley_Granger
Farley Mowat	http://en.wikipedia.org/wiki/Farley_Mowat
Faron Young	http://en.wikipedia.org/wiki/Faron_Young
Farrah Fawcett	http://en.wikipedia.org/wiki/Farrah_Fawcett
Fat Joe	http://en.wikipedia.org/wiki/Fat_Joe
Fat Mike	http://en.wikipedia.org/wiki/Fat_Mike
Fatboy Slim	http://en.wikipedia.org/wiki/Fat_Mike
Father Charles Coughlin	http://en.wikipedia.org/wiki/Father_Charles_Coughlin
Father Damien	http://en.wikipedia.org/wiki/Father_Damien
Father Joseph	http://en.wikipedia.org/wiki/Father_Joseph
Father Yod	http://en.wikipedia.org/wiki/Father_Yod
Fatmir Sejdiu	http://en.wikipedia.org/wiki/Fatmir_Sejdiu
Fats Domino	http://en.wikipedia.org/wiki/Fats_Domino
Fats Waller	http://en.wikipedia.org/wiki/Fats_Waller
Fatty Arbuckle	http://en.wikipedia.org/wiki/Fatty_Arbuckle
Faure Gnassingb�	http://en.wikipedia.org/wiki/Faure_Gnassingb%C3%A9
Faustin-Archange Touad�ra	http://en.wikipedia.org/wiki/Faustin-Archange_Touad%C3%A9ra
Fausto Vitello	http://en.wikipedia.org/wiki/Fausto_Vitello
Fawn Hall	http://en.wikipedia.org/wiki/Fawn_Hall
Fay Bainter	http://en.wikipedia.org/wiki/Fay_Bainter
Fay Vincent	http://en.wikipedia.org/wiki/Fay_Vincent
Fay Weldon	http://en.wikipedia.org/wiki/Fay_Weldon
Fay Wray	http://en.wikipedia.org/wiki/Fay_Wray
Fayard Nicholas	http://en.wikipedia.org/wiki/Fayard_Nicholas
Faye Dunaway	http://en.wikipedia.org/wiki/Faye_Dunaway
Faye Emerson	http://en.wikipedia.org/wiki/Faye_Emerson
Federico Castelluccio	http://en.wikipedia.org/wiki/Federico_Castelluccio
Federico Fellini	http://en.wikipedia.org/wiki/Federico_Fellini
Federico Garc�a Lorca	http://en.wikipedia.org/wiki/Federico_Garc%C3%ADa_Lorca
Federico Peña	http://en.wikipedia.org/wiki/Federico_Pe%C3%B1a
Fee Waybill	http://en.wikipedia.org/wiki/Fee_Waybill
Fela Kuti	http://en.wikipedia.org/wiki/Fela_Kuti
Feleti Sevele	http://en.wikipedia.org/wiki/Feleti_Sevele
Felice Cavallotti	http://en.wikipedia.org/wiki/Felice_Cavallotti
Felice Orsini	http://en.wikipedia.org/wiki/Felice_Orsini
F�licien-C�sar David	http://en.wikipedia.org/wiki/F%C3%A9licien-C%C3%A9sar_David
Felicity Huffman	http://en.wikipedia.org/wiki/Felicity_Huffman
Felicity Kendal	http://en.wikipedia.org/wiki/Felicity_Kendal
Feliks Kulov	http://en.wikipedia.org/wiki/Feliks_Kulov
Felipe Calder�n	http://en.wikipedia.org/wiki/Felipe_Calder%C3%B3n
Felisberto Hern�ndez	http://en.wikipedia.org/wiki/Felisberto_Hern%C3%A1ndez
Felix Adler	http://en.wikipedia.org/wiki/Felix_Adler_(Society_for_Ethical_Culture)
Felix Bloch	http://en.wikipedia.org/wiki/Felix_Bloch
Felix Camacho	http://en.wikipedia.org/wiki/Felix_Camacho
Felix Frankfurter	http://en.wikipedia.org/wiki/Felix_Frankfurter
Felix Mendelssohn	http://en.wikipedia.org/wiki/Felix_Mendelssohn
Felix Perez Camacho	http://en.wikipedia.org/wiki/Felix_Perez_Camacho
F�lix Rodr�guez	http://en.wikipedia.org/wiki/F%C3%A9lix_Rodr%C3%ADguez_%28Central_Intelligence_Agency%29
Felix Silla	http://en.wikipedia.org/wiki/Felix_Silla
Fenton J. A. Hort	http://en.wikipedia.org/wiki/Fenton_J._A._Hort
Ferdi Sabit Soyer	http://en.wikipedia.org/wiki/Ferdi_Sabit_Soyer
Ferdinand Braun	http://en.wikipedia.org/wiki/Ferdinand_Braun
Ferdinand Buisson	http://en.wikipedia.org/wiki/Ferdinand_Buisson
Ferdinand de Lesseps	http://en.wikipedia.org/wiki/Ferdinand_de_Lesseps
Ferdinand Foch	http://en.wikipedia.org/wiki/Ferdinand_Foch
Ferdinand Magellan	http://en.wikipedia.org/wiki/Ferdinand_Magellan
Ferdinand Marcos	http://en.wikipedia.org/wiki/Ferdinand_Marcos
Ferdinand VI	http://en.wikipedia.org/wiki/Ferdinand_VI
Ferdinand VII	http://en.wikipedia.org/wiki/Ferdinand_VII
Ferdinand von Zeppelin	http://en.wikipedia.org/wiki/Ferdinand_von_Zeppelin
Ferenc De�k	http://en.wikipedia.org/wiki/Ferenc_De%C3%A1k
Ferenc Gyurcs�ny	http://en.wikipedia.org/wiki/Ferenc_Gyurcs%C3%A1ny
Ferenc Moln�r	http://en.wikipedia.org/wiki/Ferenc_Moln%C3%A1r
Ferenc Nagy	http://en.wikipedia.org/wiki/Ferenc_Nagy
Ferenc Pusk�s	http://en.wikipedia.org/wiki/Ferenc_Pusk%C3%A1s
Fernand J. St. Germain	http://en.wikipedia.org/wiki/Fernand_J._St._Germain
Fernanda Montenegro	http://en.wikipedia.org/wiki/Fernanda_Montenegro
Fernando Alonso	http://en.wikipedia.org/wiki/Fernando_Alonso
Fernando da Piedade Dias dos Santos	http://en.wikipedia.org/wiki/Fernando_da_Piedade_Dias_dos_Santos
Fernando I	http://en.wikipedia.org/wiki/Ferdinand_I_of_Portugal
Fernando Lamas	http://en.wikipedia.org/wiki/Fernando_Lamas
Fernando Lugo	http://en.wikipedia.org/wiki/Fernando_Lugo
Fernando Pessoa	http://en.wikipedia.org/wiki/Fernando_Pessoa
Fernando Poe, Jr.	http://en.wikipedia.org/wiki/Fernando_Poe%2C_Jr.
Fernando Rey	http://en.wikipedia.org/wiki/Fernando_Rey
Fernando Valenzuela	http://en.wikipedia.org/wiki/Fernando_Valenzuela
Ferruccio Busoni	http://en.wikipedia.org/wiki/Ferruccio_Busoni
Fess Parker	http://en.wikipedia.org/wiki/Fess_Parker
Festus Mogae	http://en.wikipedia.org/wiki/Festus_Mogae
Fidel Castro	http://en.wikipedia.org/wiki/Fidel_Castro
Fidel Ramos	http://en.wikipedia.org/wiki/Fidel_Ramos
Fife Symington	http://en.wikipedia.org/wiki/Fife_Symington
Filip Vujanovic	http://en.wikipedia.org/wiki/Filip_Vujanovic
Filippo Brunelleschi	http://en.wikipedia.org/wiki/Filippo_Brunelleschi
Filoimea Telito	http://en.wikipedia.org/wiki/Filoimea_Telito
Finley Peter Dunne	http://en.wikipedia.org/wiki/Finley_Peter_Dunne
Finn Aabye	http://en.wikipedia.org/wiki/Finn_Aabye
Finola Hughes	http://en.wikipedia.org/wiki/Finola_Hughes
Fiona Apple	http://en.wikipedia.org/wiki/Fiona_Apple
Fiona Bruce	http://en.wikipedia.org/wiki/Fiona_Bruce
Fiona Mactaggart	http://en.wikipedia.org/wiki/Fiona_Mactaggart
Fiona O'Donnell	http://en.wikipedia.org/wiki/Fiona_O%27Donnell
Fiona Shaw	http://en.wikipedia.org/wiki/Fiona_Shaw
Fiorello LaGuardia	http://en.wikipedia.org/wiki/Fiorello_LaGuardia
Fisher Stevens	http://en.wikipedia.org/wiki/Fisher_Stevens
Fitz-James O'Brien	http://en.wikipedia.org/wiki/Fitz-James_O%27Brien
Flann O'Brien	http://en.wikipedia.org/wiki/Flann_O%27Brien
Flannery O'Connor	http://en.wikipedia.org/wiki/Flannery_O%27Connor
Flavius Stilicho	http://en.wikipedia.org/wiki/Flavius_Stilicho
Flavor Flav	http://en.wikipedia.org/wiki/Flavor_Flav
Flemming Ahlberg	http://en.wikipedia.org/wiki/Flemming_Ahlberg
Flip Wilson	http://en.wikipedia.org/wiki/Flip_Wilson
Flora Robson	http://en.wikipedia.org/wiki/Flora_Robson
Florence Ballard	http://en.wikipedia.org/wiki/Florence_Ballard
Florence Griffith Joyner	http://en.wikipedia.org/wiki/Florence_Griffith_Joyner
Florence Henderson	http://en.wikipedia.org/wiki/Florence_Henderson
Florence Nightingale	http://en.wikipedia.org/wiki/Florence_Nightingale
Florenz Ziegfeld	http://en.wikipedia.org/wiki/Florenz_Ziegfeld
Florian Cajori	http://en.wikipedia.org/wiki/Florian_Cajori
Florian Schneider	http://en.wikipedia.org/wiki/Florian_Schneider
Floyd Abrams	http://en.wikipedia.org/wiki/Floyd_Abrams
Floyd Cramer	http://en.wikipedia.org/wiki/Floyd_Cramer
Floyd Dell	http://en.wikipedia.org/wiki/Floyd_Dell
Floyd Patterson	http://en.wikipedia.org/wiki/Floyd_Patterson
Floyd Sneed	http://en.wikipedia.org/wiki/Floyd_Sneed
Floyd Spence	http://en.wikipedia.org/wiki/Floyd_Spence
Floyd Tillman	http://en.wikipedia.org/wiki/Floyd_Tillman
Flynt Leverett	http://en.wikipedia.org/wiki/Flynt_Leverett
Fofo I.F. Sunia	http://en.wikipedia.org/wiki/Fof%C3%B3_Iosefa_Fiti_Sunia
Ford Madox Brown	http://en.wikipedia.org/wiki/Ford_Madox_Brown
Ford Madox Ford	http://en.wikipedia.org/wiki/Ford_Madox_Ford
Ford Rainey	http://en.wikipedia.org/wiki/Ford_Rainey
Forest Whitaker	http://en.wikipedia.org/wiki/Forest_Whitaker
Forrest Tucker	http://en.wikipedia.org/wiki/Forrest_Tucker
Foster Brooks	http://en.wikipedia.org/wiki/Foster_Brooks
Fouad Siniora	http://en.wikipedia.org/wiki/Fouad_Siniora
Foxy Brown	http://en.wikipedia.org/wiki/Foxy_Brown_(singer)
Fra Angelico	http://en.wikipedia.org/wiki/Fra_Angelico
Fra Diamante	http://en.wikipedia.org/wiki/Fra_Diamante
Fra Filippo Lippi	http://en.wikipedia.org/wiki/Fra_Filippo_Lippi
Fradique de Menezes	http://en.wikipedia.org/wiki/Fradique_de_Menezes
Fran Drescher	http://en.wikipedia.org/wiki/Fran_Drescher
Fran Lebowitz	http://en.wikipedia.org/wiki/Fran_Lebowitz
Fran Tarkenton	http://en.wikipedia.org/wiki/Fran_Tarkenton
France Nuyen	http://en.wikipedia.org/wiki/France_Nuyen
Frances Bavier	http://en.wikipedia.org/wiki/Frances_Bavier
Frances Bean Cobain	http://en.wikipedia.org/wiki/Frances_Bean_Cobain
Frances Buss	http://en.wikipedia.org/wiki/Frances_Buss
Frances Conroy	http://en.wikipedia.org/wiki/Frances_Conroy
Frances Dee	http://en.wikipedia.org/wiki/Frances_Dee
Frances Drake	http://en.wikipedia.org/wiki/Frances_Drake
Frances E. W. Harper	http://en.wikipedia.org/wiki/Frances_E._W._Harper
Frances Farmer	http://en.wikipedia.org/wiki/Frances_Farmer
Frances Faye	http://en.wikipedia.org/wiki/Frances_Faye
Frances Fisher	http://en.wikipedia.org/wiki/Frances_Fisher
Frances Hodgson Burnett	http://en.wikipedia.org/wiki/Frances_Hodgson_Burnett
Frances Langford	http://en.wikipedia.org/wiki/Frances_Langford
Frances McDormand	http://en.wikipedia.org/wiki/Frances_McDormand
Frances Moore Lappe	http://en.wikipedia.org/wiki/Frances_Moore_Lappe
Frances Parkinson Keyes	http://en.wikipedia.org/wiki/Frances_Parkinson_Keyes
Frances Perkins	http://en.wikipedia.org/wiki/Frances_Perkins
Frances Rafferty	http://en.wikipedia.org/wiki/Frances_Rafferty
Frances Reid	http://en.wikipedia.org/wiki/Frances_Reid
Frances Yates	http://en.wikipedia.org/wiki/Frances_Yates
Francesca Annis	http://en.wikipedia.org/wiki/Francesca_Annis
Francesco Borromini	http://en.wikipedia.org/wiki/Francesco_Borromini
Francesco Cavalli	http://en.wikipedia.org/wiki/Francesco_Cavalli
Francesco Colonna	http://en.wikipedia.org/wiki/Francesco_Colonna
Francesco Crispi	http://en.wikipedia.org/wiki/Francesco_Crispi
Francesco Durante	http://en.wikipedia.org/wiki/Francesco_Durante
Francesco Filelfo	http://en.wikipedia.org/wiki/Francesco_Filelfo
Franchot Tone	http://en.wikipedia.org/wiki/Franchot_Tone
Francine Busby	http://en.wikipedia.org/wiki/Francine_Busby
Francis A. Walker	http://en.wikipedia.org/wiki/Francis_Amasa_Walker
Francis Arinze	http://en.wikipedia.org/wiki/Francis_Arinze
Francis Asbury	http://en.wikipedia.org/wiki/Francis_Asbury
Francis Bacon	http://en.wikipedia.org/wiki/Francis_Bacon
Francis Bacon	http://en.wikipedia.org/wiki/Francis_Bacon
Francis Baily	http://en.wikipedia.org/wiki/Francis_Baily
Francis Biddle	http://en.wikipedia.org/wiki/Francis_Biddle
Francis Crick	http://en.wikipedia.org/wiki/Francis_Crick
Francis Ford Coppola	http://en.wikipedia.org/wiki/Francis_Ford_Coppola
Francis Fukuyama	http://en.wikipedia.org/wiki/Francis_Fukuyama
Francis Galton	http://en.wikipedia.org/wiki/Francis_Galton
Francis Gary Powers	http://en.wikipedia.org/wiki/Francis_Gary_Powers
Francis Healy	http://en.wikipedia.org/wiki/Francis_Healy
Francis Henry Underwood	http://en.wikipedia.org/wiki/Francis_Henry_Underwood
Francis Hopkinson	http://en.wikipedia.org/wiki/Francis_Hopkinson
Francis Horner	http://en.wikipedia.org/wiki/Francis_Horner
Francis I	http://en.wikipedia.org/wiki/Francis_I_of_France
Francis II	http://en.wikipedia.org/wiki/Francis_II_of_France
Francis Ledwidge	http://en.wikipedia.org/wiki/Francis_Ledwidge
Francis Lewis	http://en.wikipedia.org/wiki/Francis_Lewis
Francis Marion	http://en.wikipedia.org/wiki/Francis_Marion
Francis Maude	http://en.wikipedia.org/wiki/Francis_Maude
Francis Parkman	http://en.wikipedia.org/wiki/Francis_Parkman
Francis Poulenc	http://en.wikipedia.org/wiki/Francis_Poulenc
Francis Rawdon-Hastings	http://en.wikipedia.org/wiki/Francis_Rawdon-Hastings
Francis Scott Key	http://en.wikipedia.org/wiki/Francis_Scott_Key
Francis Steegmuller	http://en.wikipedia.org/wiki/Francis_Steegmuller
Francis Turner Palgrave	http://en.wikipedia.org/wiki/Francis_Turner_Palgrave
Francis W. Aston	http://en.wikipedia.org/wiki/Francis_W._Aston
Francis X. Bushman	http://en.wikipedia.org/wiki/Francis_X._Bushman
Francisco de Goya	http://en.wikipedia.org/wiki/Francisco_de_Goya
Francisco Franco	http://en.wikipedia.org/wiki/Francisco_Franco
Francisco Jim�nez de Cisneros	http://en.wikipedia.org/wiki/Francisco_Jim%C3%A9nez_de_Cisneros
Francisco Pizarro	http://en.wikipedia.org/wiki/Francisco_Pizarro
Francisco Su�rez	http://en.wikipedia.org/wiki/Francisco_Su%C3%A1rez
Francisco V�squez de Coronado	http://en.wikipedia.org/wiki/Francisco_V%C3%A1zquez_de_Coronado
Francisco Zurbar�n	http://en.wikipedia.org/wiki/Francisco_de_Zurbar%C3%A1n
Franco Ambrosetti	http://en.wikipedia.org/wiki/Franco_Ambrosetti
Franco Harris	http://en.wikipedia.org/wiki/Franco_Harris
Franco Nero	http://en.wikipedia.org/wiki/Franco_Nero
Franco Zeffirelli	http://en.wikipedia.org/wiki/Franco_Zeffirelli
Fran�ois Arago	http://en.wikipedia.org/wiki/Fran%C3%A7ois_Arago
Francois Bozize	http://en.wikipedia.org/wiki/Francois_Bozize
Fran�ois Boziz�	http://en.wikipedia.org/wiki/Fran%C3%A7ois_Boziz%C3%A9
Fran�ois Couperin	http://en.wikipedia.org/wiki/Fran%C3%A7ois_Couperin
Fran�ois de la Rochefoucauld	http://en.wikipedia.org/wiki/Fran%C3%A7ois_de_la_Rochefoucauld
Fran�ois de Malherbe	http://en.wikipedia.org/wiki/Fran%C3%A7ois_de_Malherbe
Fran�ois Duvalier	http://en.wikipedia.org/wiki/Fran%C3%A7ois_Duvalier
Fran�ois F�nelon	http://en.wikipedia.org/wiki/Fran%C3%A7ois_F%C3%A9nelon
Fran�ois Fillon	http://en.wikipedia.org/wiki/Fran%C3%A7ois_Fillon
Fran�ois Girardon	http://en.wikipedia.org/wiki/Fran%C3%A7ois_Girardon
Fran�ois Guizot	http://en.wikipedia.org/wiki/Fran%C3%A7ois_Guizot
Fran�ois Hanriot	http://en.wikipedia.org/wiki/Fran%C3%A7ois_Hanriot
Fran�ois Hotman	http://en.wikipedia.org/wiki/Fran%C3%A7ois_Hotman
Fran�ois Mansart	http://en.wikipedia.org/wiki/Fran%C3%A7ois_Mansart
Fran�ois Mauriac	http://en.wikipedia.org/wiki/Fran%C3%A7ois_Mauriac
Fran�ois Mitterrand	http://en.wikipedia.org/wiki/Fran%C3%A7ois_Mitterrand
Fran�ois Rabelais	http://en.wikipedia.org/wiki/Fran%C3%A7ois_Rabelais
Fran�ois Truffaut	http://en.wikipedia.org/wiki/Fran%C3%A7ois_Truffaut
Fran�oise Hardy	http://en.wikipedia.org/wiki/Fran%C3%A7oise_Hardy
Fran�ois-Ren� de Chateaubriand	http://en.wikipedia.org/wiki/Fran%C3%A7ois-Ren%C3%A9_de_Chateaubriand
Franjo Tudjman	http://en.wikipedia.org/wiki/Franjo_Tudjman
Frank Abney Hastings	http://en.wikipedia.org/wiki/Frank_Abney_Hastings
Frank Adonis	http://en.wikipedia.org/wiki/Frank_Adonis
Frank Agrama	http://en.wikipedia.org/wiki/Frank_Agrama
Frank Annunzio	http://en.wikipedia.org/wiki/Frank_Annunzio
Frank B. Kellogg	http://en.wikipedia.org/wiki/Frank_B._Kellogg
Frank B. Morrison	http://en.wikipedia.org/wiki/Frank_B._Morrison
Frank Bainimarama	http://en.wikipedia.org/wiki/Frank_Bainimarama
Frank Ballance	http://en.wikipedia.org/wiki/Frank_Ballance
Frank Bidart	http://en.wikipedia.org/wiki/Frank_Bidart
Frank Biondi	http://en.wikipedia.org/wiki/Frank_Biondi
Frank Black	http://en.wikipedia.org/wiki/Frank_Black
Frank Bonner	http://en.wikipedia.org/wiki/Frank_Bonner
Frank Borman	http://en.wikipedia.org/wiki/Frank_Borman
Frank Borzage	http://en.wikipedia.org/wiki/Frank_Borzage
Frank Bruni	http://en.wikipedia.org/wiki/Frank_Bruni
Frank Cady	http://en.wikipedia.org/wiki/Frank_Cady
Frank Capra	http://en.wikipedia.org/wiki/Frank_Capra
Frank Carlucci	http://en.wikipedia.org/wiki/Frank_Carlucci
Frank Carson	http://en.wikipedia.org/wiki/Frank_Carson
Frank Church	http://en.wikipedia.org/wiki/Frank_Church
Frank Corder	http://en.wikipedia.org/wiki/Frank_Eugene_Corder
Frank Darabont	http://en.wikipedia.org/wiki/Frank_Darabont
Frank De Vol	http://en.wikipedia.org/wiki/Frank_De_Vol
Frank DeKova	http://en.wikipedia.org/wiki/Frank_DeKova
Frank Dobson	http://en.wikipedia.org/wiki/Frank_Dobson
Frank Doran	http://en.wikipedia.org/wiki/Frank_Doran_(UK_politician)
Frank Doubleday	http://en.wikipedia.org/wiki/Frank_Doubleday
Frank Farian	http://en.wikipedia.org/wiki/Frank_Farian
Frank Field	http://en.wikipedia.org/wiki/Frank_Field_(politician)
Frank Frazetta	http://en.wikipedia.org/wiki/Frank_Frazetta
Frank G. Clement	http://en.wikipedia.org/wiki/Frank_G._Clement
Frank Gaffney	http://en.wikipedia.org/wiki/Frank_Gaffney
Frank Gannett	http://en.wikipedia.org/wiki/Frank_Gannett
Frank Gehry	http://en.wikipedia.org/wiki/Frank_Gehry
Frank Gifford	http://en.wikipedia.org/wiki/Frank_Gifford
Frank Gorshin	http://en.wikipedia.org/wiki/Frank_Gorshin
Frank H. Murkowski	http://en.wikipedia.org/wiki/Frank_H._Murkowski
Frank Harris	http://en.wikipedia.org/wiki/Frank_Harris
Frank Herbert	http://en.wikipedia.org/wiki/Frank_Herbert
Frank Horton	http://en.wikipedia.org/wiki/Frank_Horton
Frank Hsieh	http://en.wikipedia.org/wiki/Frank_Hsieh
Frank Iero	http://en.wikipedia.org/wiki/Frank_Iero
Frank Jordan	http://en.wikipedia.org/wiki/Frank_Jordan
Frank Kelly Freas	http://en.wikipedia.org/wiki/Frank_Kelly_Freas
Frank Kermode	http://en.wikipedia.org/wiki/Frank_Kermode
Frank King	http://en.wikipedia.org/wiki/Frank_King_(cartoonist)
Frank Kratovil	http://en.wikipedia.org/wiki/Frank_Kratovil
Frank Lampard	http://en.wikipedia.org/wiki/Frank_Lampard
Frank Langella	http://en.wikipedia.org/wiki/Frank_Langella
Frank Lautenberg	http://en.wikipedia.org/wiki/Frank_Lautenberg
Frank Lloyd	http://en.wikipedia.org/wiki/Frank_Lloyd
Frank Lloyd Wright	http://en.wikipedia.org/wiki/Frank_Lloyd_Wright
Frank LoBiondo	http://en.wikipedia.org/wiki/Frank_LoBiondo
Frank Lorenzo	http://en.wikipedia.org/wiki/Frank_Lorenzo
Frank Lucas	http://en.wikipedia.org/wiki/Frank_Lucas_(politician)
Frank Luntz	http://en.wikipedia.org/wiki/Frank_Luntz
Frank McCloskey	http://en.wikipedia.org/wiki/Frank_McCloskey
Frank McCourt	http://en.wikipedia.org/wiki/Frank_McCourt
Frank Miller	http://en.wikipedia.org/wiki/Frank_Miller_(comics)
Frank Morgan	http://en.wikipedia.org/wiki/Frank_Morgan
Frank Murkowski	http://en.wikipedia.org/wiki/Frank_Murkowski
Frank Murkowski	http://en.wikipedia.org/wiki/Frank_Murkowski
Frank Norris	http://en.wikipedia.org/wiki/Frank_Norris
Frank O'Connor	http://en.wikipedia.org/wiki/Frank_O%27Connor
Frank O'Hara	http://en.wikipedia.org/wiki/Frank_O%27Hara
Frank Oppenheimer	http://en.wikipedia.org/wiki/Frank_Oppenheimer
Frank Oz	http://en.wikipedia.org/wiki/Frank_Oz
Frank Pallone	http://en.wikipedia.org/wiki/Frank_Pallone
Frank Perdue	http://en.wikipedia.org/wiki/Frank_Perdue
Frank Quattrone	http://en.wikipedia.org/wiki/Frank_Quattrone
Frank R. Lautenberg	http://en.wikipedia.org/wiki/Frank_R._Lautenberg
Frank R. Wolf	http://en.wikipedia.org/wiki/Frank_R._Wolf
Frank Reynolds	http://en.wikipedia.org/wiki/Frank_Reynolds
Frank Rich	http://en.wikipedia.org/wiki/Frank_Rich
Frank Robinson	http://en.wikipedia.org/wiki/Frank_Robinson
Frank Rosolino	http://en.wikipedia.org/wiki/Frank_Rosolino
Frank Roy	http://en.wikipedia.org/wiki/Frank_Roy
Frank Serpico	http://en.wikipedia.org/wiki/Frank_Serpico
Frank Sesno	http://en.wikipedia.org/wiki/Frank_Sesno
Frank Shakespeare	http://en.wikipedia.org/wiki/Frank_Shakespeare
Frank Sinatra	http://en.wikipedia.org/wiki/Frank_Sinatra
Frank Sinatra, Jr.	http://en.wikipedia.org/wiki/Frank_Sinatra%2C_Jr.
Frank Stallone	http://en.wikipedia.org/wiki/Frank_Stallone
Frank Sutton	http://en.wikipedia.org/wiki/Frank_Sutton
Frank Tashlin	http://en.wikipedia.org/wiki/Frank_Tashlin
Frank Turner	http://en.wikipedia.org/wiki/Frank_Turner
Frank Walker	http://en.wikipedia.org/wiki/Frank_Walker_(Jersey_politician)
Frank Wedekind	http://en.wikipedia.org/wiki/Frank_Wedekind
Frank Whaley	http://en.wikipedia.org/wiki/Frank_Whaley
Frank Wolf	http://en.wikipedia.org/wiki/Frank_Wolf
Frank Yerby	http://en.wikipedia.org/wiki/Frank_Yerby
Frank Zappa	http://en.wikipedia.org/wiki/Frank_Zappa
Frankie Avalon	http://en.wikipedia.org/wiki/Frankie_Avalon
Frankie Darro	http://en.wikipedia.org/wiki/Frankie_Darro
Frankie Faison	http://en.wikipedia.org/wiki/Frankie_Faison
Frankie Frisch	http://en.wikipedia.org/wiki/Frankie_Frisch
Frankie Howerd	http://en.wikipedia.org/wiki/Frankie_Howerd
Frankie J	http://en.wikipedia.org/wiki/Frankie_J
Frankie Laine	http://en.wikipedia.org/wiki/Frankie_Laine
Frankie Lymon	http://en.wikipedia.org/wiki/Frankie_Lymon
Frankie Muniz	http://en.wikipedia.org/wiki/Frankie_Mu%C3%B1iz
Frankie Valli	http://en.wikipedia.org/wiki/Frankie_Valli
Frankie Yankovic	http://en.wikipedia.org/wiki/Frankie_Yankovic
Franklin Adreon	http://en.wikipedia.org/wiki/Franklin_Adreon
Franklin Cover	http://en.wikipedia.org/wiki/Franklin_Cover
Franklin D. Roosevelt	http://en.wikipedia.org/wiki/Franklin_D._Roosevelt
Franklin J. Schaffner	http://en.wikipedia.org/wiki/Franklin_J._Schaffner
Franklin K. Lane	http://en.wikipedia.org/wiki/Franklin_K._Lane
Franklin Pierce	http://en.wikipedia.org/wiki/Franklin_Pierce
Franklin Pierce Adams	http://en.wikipedia.org/wiki/Franklin_Pierce_Adams
Franklin Raines	http://en.wikipedia.org/wiki/Franklin_Raines
Frans Hals	http://en.wikipedia.org/wiki/Frans_Hals
Franz Aigner	http://en.wikipedia.org/wiki/Franz_Aigner_%28footballer%29
Franz Anton Mesmer	http://en.wikipedia.org/wiki/Franz_Anton_Mesmer
Franz Beckenbauer	http://en.wikipedia.org/wiki/Franz_Beckenbauer
Franz Boas	http://en.wikipedia.org/wiki/Franz_Boas
Franz Bopp	http://en.wikipedia.org/wiki/Franz_Bopp
Franz Ferdinand	http://en.wikipedia.org/wiki/Franz_Ferdinand
Franz Grillparzer	http://en.wikipedia.org/wiki/Franz_Grillparzer
Franz Guertner	http://en.wikipedia.org/wiki/Franz_Guertner
Franz Halder	http://en.wikipedia.org/wiki/Franz_Halder
Franz Joseph Gall	http://en.wikipedia.org/wiki/Franz_Joseph_Gall
Franz Kafka	http://en.wikipedia.org/wiki/Franz_Kafka
Franz Kline	http://en.wikipedia.org/wiki/Franz_Kline
Franz Kotzwara	http://en.wikipedia.org/wiki/Franz_Kotzwara
Franz Liszt	http://en.wikipedia.org/wiki/Franz_Liszt
Franz M�ntefering	http://en.wikipedia.org/wiki/Franz_M%C3%Bcntefering
Franz Ritter von Hauer	http://en.wikipedia.org/wiki/Franz_Ritter_von_Hauer
Franz Schubert	http://en.wikipedia.org/wiki/Franz_Schubert
Franz von Papen	http://en.wikipedia.org/wiki/Franz_von_Papen
Franz Vranitzky	http://en.wikipedia.org/wiki/Franz_Vranitzky
Franz Waxman	http://en.wikipedia.org/wiki/Franz_Waxman
Fred A. Seaton	http://en.wikipedia.org/wiki/Fred_A._Seaton
Fred Allen	http://en.wikipedia.org/wiki/Fred_Allen
Fred Armisen	http://en.wikipedia.org/wiki/Fred_Armisen
Fred Astaire	http://en.wikipedia.org/wiki/Fred_Astaire
Fred Barnes	http://en.wikipedia.org/wiki/Fred_Barnes_(journalist)
Fred Berry	http://en.wikipedia.org/wiki/Fred_Berry
Fred Bodsworth	http://en.wikipedia.org/wiki/Fred_Bodsworth
Fred Brooks	http://en.wikipedia.org/wiki/Fred_Brooks
Fred C. Koch	http://en.wikipedia.org/wiki/Fred_C._Koch
Fred Couples	http://en.wikipedia.org/wiki/Fred_Couples
Fred Dryer	http://en.wikipedia.org/wiki/Fred_Dryer
Fred Durst	http://en.wikipedia.org/wiki/Fred_Durst
Fred Ebb	http://en.wikipedia.org/wiki/Fred_Ebb
Fred F. Fielding	http://en.wikipedia.org/wiki/Fred_F._Fielding
Fred Friendly	http://en.wikipedia.org/wiki/Fred_Friendly
Fred Frith	http://en.wikipedia.org/wiki/Fred_Frith
Fred Grandy	http://en.wikipedia.org/wiki/Fred_Grandy
Fred Gwynne	http://en.wikipedia.org/wiki/Fred_Gwynne
Fred Hoyle	http://en.wikipedia.org/wiki/Fred_Hoyle
Fred J. Eckert	http://en.wikipedia.org/wiki/Fred_J._Eckert
Fred Karlin	http://en.wikipedia.org/wiki/Fred_Karlin
Fred LaRue	http://en.wikipedia.org/wiki/Fred_LaRue
Fred Leuchter, Jr.	http://en.wikipedia.org/wiki/Fred_A._Leuchter
Fred MacMurray	http://en.wikipedia.org/wiki/Fred_MacMurray
Fred Malek	http://en.wikipedia.org/wiki/Fred_Malek
Fred Phelps	http://en.wikipedia.org/wiki/Fred_Phelps
Fred Quimby	http://en.wikipedia.org/wiki/Fred_Quimby
Fred Rogers	http://en.wikipedia.org/wiki/Fred_Rogers
Fred Rogers	http://en.wikipedia.org/wiki/Fred_Rogers
Fred Saberhagen	http://en.wikipedia.org/wiki/Fred_Saberhagen
Fred Savage	http://en.wikipedia.org/wiki/Fred_Savage
Fred Schepisi	http://en.wikipedia.org/wiki/Fred_Schepisi
Fred Schneider	http://en.wikipedia.org/wiki/Fred_Schneider
Fred Silverman	http://en.wikipedia.org/wiki/Fred_Silverman
Fred Thompson	http://en.wikipedia.org/wiki/Fred_Thompson
Fred Turner	http://en.wikipedia.org/wiki/Fred_Turner_(musician)
Fred Upton	http://en.wikipedia.org/wiki/Fred_Upton
Fred Vinson	http://en.wikipedia.org/wiki/Fred_M._Vinson
Fred Ward	http://en.wikipedia.org/wiki/Fred_Ward
Fred Waring	http://en.wikipedia.org/wiki/Fred_Waring
Fred Whipple	http://en.wikipedia.org/wiki/Fred_Whipple
Fred Willard	http://en.wikipedia.org/wiki/Fred_Willard
Fred Williamson	http://en.wikipedia.org/wiki/Fred_Williamson
Fred Zinnemann	http://en.wikipedia.org/wiki/Fred_Zinnemann
Freddie Bartholomew	http://en.wikipedia.org/wiki/Freddie_Bartholomew
Freddie Hubbard	http://en.wikipedia.org/wiki/Freddie_Hubbard
Freddie Jackson	http://en.wikipedia.org/wiki/Freddie_Jackson
Freddie Laker	http://en.wikipedia.org/wiki/Freddie_Laker
Freddie Mercury	http://en.wikipedia.org/wiki/Freddie_Mercury
Freddie Prinze	http://en.wikipedia.org/wiki/Freddie_Prinze
Freddie Prinze, Jr.	http://en.wikipedia.org/wiki/Freddie_Prinze%2C_Jr.
Freddie Young	http://en.wikipedia.org/wiki/Freddie_Young
Freddy Fender	http://en.wikipedia.org/wiki/Freddy_Fender
Frederic Chopin	http://en.wikipedia.org/wiki/Frederic_Chopin
Frederic Jameson	http://en.wikipedia.org/wiki/Frederic_Jameson
Fr�d�ric Joliot	http://en.wikipedia.org/wiki/Fr%C3%A9d%C3%A9ric_Joliot
Frederic Manning	http://en.wikipedia.org/wiki/Frederic_Manning
Fr�d�ric Mistral	http://en.wikipedia.org/wiki/Fr%C3%A9d%C3%A9ric_Mistral
Fr�d�ric Passy	http://en.wikipedia.org/wiki/Fr%C3%A9d%C3%A9ric_Passy
Frederic Prokosch	http://en.wikipedia.org/wiki/Frederic_Prokosch
Frederic Remington	http://en.wikipedia.org/wiki/Frederic_Remington
Frederic W. Goudy	http://en.wikipedia.org/wiki/Frederic_W._Goudy
Frederick Barthelme	http://en.wikipedia.org/wiki/Frederick_Barthelme
Frederick Buechner	http://en.wikipedia.org/wiki/Frederick_Buechner
Frederick Busch	http://en.wikipedia.org/wiki/Frederick_Busch
Frederick De Cordova	http://en.wikipedia.org/wiki/Frederick_De_Cordova
Frederick Delius	http://en.wikipedia.org/wiki/Frederick_Delius
Frederick Denison Maurice	http://en.wikipedia.org/wiki/Frederick_Denison_Maurice
Frederick Douglass	http://en.wikipedia.org/wiki/Frederick_Douglass
Frederick Forsyth	http://en.wikipedia.org/wiki/Frederick_Forsyth
Frederick Goodwin	http://en.wikipedia.org/wiki/Frederick_Tutu_Goodwin
Frederick Jackson Turner	http://en.wikipedia.org/wiki/Frederick_Jackson_Turner
Frederick K. C. Price	http://en.wikipedia.org/wiki/Frederick_Jackson_Turner
Frederick Law Olmsted	http://en.wikipedia.org/wiki/Frederick_Law_Olmsted
Frederick Leighton	http://en.wikipedia.org/wiki/Frederick_Leighton
Frederick Lewis Allen	http://en.wikipedia.org/wiki/Frederick_Lewis_Allen
Frederick Lonsdale	http://en.wikipedia.org/wiki/Frederick_Lonsdale
Frederick Reines	http://en.wikipedia.org/wiki/Frederick_Reines
Frederick Ryan, Jr.	http://en.wikipedia.org/wiki/Fred_Ryan
Frederick Sanger	http://en.wikipedia.org/wiki/Frederick_Sanger
Frederick Soddy	http://en.wikipedia.org/wiki/Frederick_Soddy
Frederick Temple	http://en.wikipedia.org/wiki/Frederick_Temple
Frederick the Great	http://en.wikipedia.org/wiki/Frederick_the_Great
Frederick The Wise	http://en.wikipedia.org/wiki/Frederick_The_Wise
Frederik Pohl	http://en.wikipedia.org/wiki/Frederik_Pohl
Fredis Refunjol	http://en.wikipedia.org/wiki/Fredis_Refunjol
Fredric March	http://en.wikipedia.org/wiki/Fredric_March
Fredrik Bajer	http://en.wikipedia.org/wiki/Fredrik_Bajer
Fredrik Reinfeldt	http://en.wikipedia.org/wiki/Fredrik_Reinfeldt
Freeman Dyson	http://en.wikipedia.org/wiki/Freeman_Dyson
French Stewart	http://en.wikipedia.org/wiki/French_Stewart
Frenchie Davis	http://en.wikipedia.org/wiki/Frenchie_Davis
Frida Kahlo	http://en.wikipedia.org/wiki/Frida_Kahlo
Fridtjof Nansen	http://en.wikipedia.org/wiki/Fridtjof_Nansen
Friederich Konrad Hornemann	http://en.wikipedia.org/wiki/Friederich_Konrad_Hornemann
Friedrich August Kekul�	http://en.wikipedia.org/wiki/Friedrich_August_Kekul%C3%A9
Friedrich Bergius	http://en.wikipedia.org/wiki/Friedrich_Bergius
Friedrich Ebert	http://en.wikipedia.org/wiki/Friedrich_Ebert
Friedrich Engels	http://en.wikipedia.org/wiki/Friedrich_Engels
Friedrich Georg Wilhelm Struve	http://en.wikipedia.org/wiki/Friedrich_Georg_Wilhelm_Struve
Friedrich Gottlieb Klopstock	http://en.wikipedia.org/wiki/Friedrich_Gottlieb_Klopstock
Friedrich Hebbel	http://en.wikipedia.org/wiki/Friedrich_Hebbel
Friedrich Heinrich Jacobi	http://en.wikipedia.org/wiki/Friedrich_Heinrich_Jacobi
Friedrich H�lderlin	http://en.wikipedia.org/wiki/Friedrich_H%C3%B6lderlin
Friedrich Hund	http://en.wikipedia.org/wiki/Friedrich_Hund
Friedrich Leibacher	http://en.wikipedia.org/wiki/Friedrich_Leibacher
Friedrich Maximilian Klinger	http://en.wikipedia.org/wiki/Friedrich_Maximilian_Klinger
Friedrich Merz	http://en.wikipedia.org/wiki/Friedrich_Merz
Friedrich Myconius	http://en.wikipedia.org/wiki/Friedrich_Myconius
Friedrich Nietzsche	http://en.wikipedia.org/wiki/Friedrich_Nietzsche
Friedrich Olbricht	http://en.wikipedia.org/wiki/Friedrich_Olbricht
Friedrich Paulus	http://en.wikipedia.org/wiki/Friedrich_Paulus
Friedrich Schleiermacher	http://en.wikipedia.org/wiki/Friedrich_Schleiermacher
Friedrich von Hagedorn	http://en.wikipedia.org/wiki/Friedrich_von_Hagedorn
Friedrich von Holstein	http://en.wikipedia.org/wiki/Friedrich_von_Holstein
Friedrich von Schiller	http://en.wikipedia.org/wiki/Friedrich_von_Schiller
Friedrich von Schlegel	http://en.wikipedia.org/wiki/Friedrich_von_Schlegel
Friedrich Wilhelm August Argelander	http://en.wikipedia.org/wiki/Friedrich_Wilhelm_August_Argelander
Friedrich Wilhelm Bessel	http://en.wikipedia.org/wiki/Friedrich_Wilhelm_Bessel
Friedrich Wilhelm Joseph von Schelling	http://en.wikipedia.org/wiki/Friedrich_Wilhelm_Joseph_von_Schelling
Friedrich W�hler	http://en.wikipedia.org/wiki/Friedrich_W%C3%B6hler
Frits Goedgedrag	http://en.wikipedia.org/wiki/Frits_Goedgedrag
Frits Zernike	http://en.wikipedia.org/wiki/Frits_Zernike
Fritz Albrecht	http://en.wikipedia.org/wiki/Fritz_Albrecht
Fritz Feld	http://en.wikipedia.org/wiki/Fritz_Feld
Fritz Haber	http://en.wikipedia.org/wiki/Fritz_Haber
Fritz Hollings	http://en.wikipedia.org/wiki/Fritz_Hollings
Fritz Kolbe	http://en.wikipedia.org/wiki/Fritz_Kolbe
Fritz Lang	http://en.wikipedia.org/wiki/Fritz_Lang
Fritz Leiber	http://en.wikipedia.org/wiki/Fritz_Leiber
Fritz Pregl	http://en.wikipedia.org/wiki/Fritz_Pregl
Fritz Sauckel	http://en.wikipedia.org/wiki/Fritz_Sauckel
Fritz Todt	http://en.wikipedia.org/wiki/Fritz_Todt
Fritz Weaver	http://en.wikipedia.org/wiki/Fritz_Weaver
Friz Freleng	http://en.wikipedia.org/wiki/Friz_Freleng
Fromental Hal�vy	http://en.wikipedia.org/wiki/Fromental_Hal%C3%A9vy
Fulgencio Batista	http://en.wikipedia.org/wiki/Fulgencio_Batista
Fulke Greville	http://en.wikipedia.org/wiki/Fulke_Greville
Fuzzy Zoeller	http://en.wikipedia.org/wiki/Fuzzy_Zoeller
Fyodor Dostoevsky	http://en.wikipedia.org/wiki/Fyodor_Dostoevsky
Fyodor Tyutchev	http://en.wikipedia.org/wiki/Fyodor_Tyutchev
Fyvush Finkel	http://en.wikipedia.org/wiki/Fyvush_Finkel
G. E. Moore	http://en.wikipedia.org/wiki/G._E._Moore
G. E. Smith	http://en.wikipedia.org/wiki/G._E._Smith
G. G. Allin	http://en.wikipedia.org/wiki/G._G._Allin
G. Gordon Liddy	http://en.wikipedia.org/wiki/G._Gordon_Liddy
G. Gordon Liddy	http://en.wikipedia.org/wiki/G._Gordon_Liddy
G. I. Gurdjieff	http://en.wikipedia.org/wiki/G._I._Gurdjieff
G. K. Chesterton	http://en.wikipedia.org/wiki/G._K._Chesterton
G. M. Trevelyan	http://en.wikipedia.org/wiki/G._M._Trevelyan
G. W. Bailey	http://en.wikipedia.org/wiki/G._W._Bailey
G. W. Bitzer	http://en.wikipedia.org/wiki/G._W._Bitzer
G. William Whitehurst	http://en.wikipedia.org/wiki/G._William_Whitehurst
G.V. Montgomery	http://en.wikipedia.org/wiki/G.V._Montgomery
Gabby Hayes	http://en.wikipedia.org/wiki/Gabby_Hayes
Gabe Kaplan	http://en.wikipedia.org/wiki/Gabe_Kaplan
Gabor Szabo	http://en.wikipedia.org/wiki/Gabor_Szabo
Gabriel Alonso de Herrera	http://en.wikipedia.org/wiki/Gabriel_Alonso_de_Herrera
Gabriel Byrne	http://en.wikipedia.org/wiki/Gabriel_Byrne
Gabriel Daniel Fahrenheit	http://en.wikipedia.org/wiki/Gabriel_Daniel_Fahrenheit
Gabriel Faur�	http://en.wikipedia.org/wiki/Gabriel_Faur%C3%A9
Gabriel Garc�a M�rquez	http://en.wikipedia.org/wiki/Gabriel_Garc%C3%ADa_M%C3%A1rquez
Gabriel Harvey	http://en.wikipedia.org/wiki/Gabriel_Harvey
Gabriel Lippmann	http://en.wikipedia.org/wiki/Gabriel_Lippmann
Gabriel Tarde	http://en.wikipedia.org/wiki/Gabriel_Tarde
Gabriela Mistral	http://en.wikipedia.org/wiki/Gabriela_Mistral
Gabriele D'Annunzio	http://en.wikipedia.org/wiki/Gabriele_D%27Annunzio
Gabriele Falloppio	http://en.wikipedia.org/wiki/Gabriele_Falloppio
Gabrielle Anwar	http://en.wikipedia.org/wiki/Gabrielle_Anwar
Gabrielle Giffords	http://en.wikipedia.org/wiki/Gabrielle_Giffords
Gabrielle Union	http://en.wikipedia.org/wiki/Gabrielle_Union
Gaby Hoffmann	http://en.wikipedia.org/wiki/Gaby_Hoffmann
Gael Garc�a Bernal	http://en.wikipedia.org/wiki/Gael_Garc%C3%ADa_Bernal
Gaetano Badalamenti	http://en.wikipedia.org/wiki/Gaetano_Badalamenti
Gaetano Donizetti	http://en.wikipedia.org/wiki/Gaetano_Donizetti
Gail Ann Dorsey	http://en.wikipedia.org/wiki/Gail_Ann_Dorsey
Gail O'Grady	http://en.wikipedia.org/wiki/Gail_O%27Grady
Gail Russell	http://en.wikipedia.org/wiki/Gail_Russell
Gaius Lucilius	http://en.wikipedia.org/wiki/Gaius_Lucilius
Gaius Marius	http://en.wikipedia.org/wiki/Gaius_Marius
Gale A. Norton	http://en.wikipedia.org/wiki/Gale_A._Norton
Gale Gordon	http://en.wikipedia.org/wiki/Gale_Gordon
Gale Harold	http://en.wikipedia.org/wiki/Gale_Harold
Gale Sondergaard	http://en.wikipedia.org/wiki/Gale_Sondergaard
Gale Storm	http://en.wikipedia.org/wiki/Gale_Storm
Galileo Ferraris	http://en.wikipedia.org/wiki/Galileo_Ferraris
Galileo Galilei	http://en.wikipedia.org/wiki/Galileo_Galilei
Galway Kinnell	http://en.wikipedia.org/wiki/Galway_Kinnell
Gamal Abdel-Nasser	http://en.wikipedia.org/wiki/Gamal_Abdel-Nasser
Gamaliel Bailey	http://en.wikipedia.org/wiki/Gamaliel_Bailey
Gao Xingjian	http://en.wikipedia.org/wiki/Gao_Xingjian
Gareth Johnson	http://en.wikipedia.org/wiki/Gareth_Johnson
Gareth Thomas	http://en.wikipedia.org/wiki/Gareth_Thomas_(English_politician)
Garfield Sobers	http://en.wikipedia.org/wiki/Garfield_Sobers
Garnet Mimms	http://en.wikipedia.org/wiki/Garnet_Mimms
Garret A. Hobart	http://en.wikipedia.org/wiki/Garret_A._Hobart
Garret FitzGerald	http://en.wikipedia.org/wiki/Garret_FitzGerald
Garrett Morris	http://en.wikipedia.org/wiki/Garrett_Morris
Garrison Keillor	http://en.wikipedia.org/wiki/Garrison_Keillor
Garry Cobain	http://en.wikipedia.org/wiki/Garry_Cobain
Garry Kasparov	http://en.wikipedia.org/wiki/Garry_Kasparov
Garry Marshall	http://en.wikipedia.org/wiki/Garry_Marshall
Garry Shandling	http://en.wikipedia.org/wiki/Garry_Shandling
Garry Trudeau	http://en.wikipedia.org/wiki/Garry_Trudeau
Garry Wills	http://en.wikipedia.org/wiki/Garry_Wills
Garson Kanin	http://en.wikipedia.org/wiki/Garson_Kanin
Garth Brooks	http://en.wikipedia.org/wiki/Garth_Brooks
Garth Ennis	http://en.wikipedia.org/wiki/Garth_Ennis
Garth Hudson	http://en.wikipedia.org/wiki/Garth_Hudson
Gary "U.S." Bonds	http://en.wikipedia.org/wiki/Gary_%22U.S.%22_Bonds
Gary Ackerman	http://en.wikipedia.org/wiki/Gary_Ackerman
Gary Aldrich	http://en.wikipedia.org/wiki/Gary_Aldrich
Gary Anthony Williams	http://en.wikipedia.org/wiki/Gary_Anthony_Williams
Gary Bauer	http://en.wikipedia.org/wiki/Gary_Bauer
Gary Burghoff	http://en.wikipedia.org/wiki/Gary_Burghoff
Gary Burton	http://en.wikipedia.org/wiki/Gary_Burton
Gary Busey	http://en.wikipedia.org/wiki/Gary_Busey
Gary Cherone	http://en.wikipedia.org/wiki/Gary_Cherone
Gary Cole	http://en.wikipedia.org/wiki/Gary_Cole
Gary Coleman	http://en.wikipedia.org/wiki/Gary_Coleman
Gary Collins	http://en.wikipedia.org/wiki/Gary_Collins_(actor)
Gary Condit	http://en.wikipedia.org/wiki/Gary_Condit
Gary Cooper	http://en.wikipedia.org/wiki/Gary_Cooper
Gary Crosby	http://en.wikipedia.org/wiki/Gary_Crosby_(actor)
Gary Dell'Abate	http://en.wikipedia.org/wiki/Gary_Dell%27Abate
Gary Dourdan	http://en.wikipedia.org/wiki/Gary_Dourdan
Gary Gilmore	http://en.wikipedia.org/wiki/Gary_Gilmore
Gary Glitter	http://en.wikipedia.org/wiki/Gary_Glitter
Gary Gygax	http://en.wikipedia.org/wiki/Gary_Gygax
Gary Hart	http://en.wikipedia.org/wiki/Gary_Hart
Gary Hart	http://en.wikipedia.org/wiki/Gary_Hart
Gary Hirte	http://en.wikipedia.org/wiki/Murder_of_Glenn_Kopitske
Gary Kildall	http://en.wikipedia.org/wiki/Gary_Kildall
Gary L. Ackerman	http://en.wikipedia.org/wiki/Gary_L._Ackerman
Gary Langan	http://en.wikipedia.org/wiki/Gary_Langan
Gary Larson	http://en.wikipedia.org/wiki/Gary_Larson
Gary Leon Ridgway	http://en.wikipedia.org/wiki/Gary_Leon_Ridgway
Gary Lineker	http://en.wikipedia.org/wiki/Gary_Lineker
Gary Locke	http://en.wikipedia.org/wiki/Gary_Locke
Gary Lockwood	http://en.wikipedia.org/wiki/Gary_Lockwood
Gary Lucas	http://en.wikipedia.org/wiki/Gary_Lucas
Gary Miller	http://en.wikipedia.org/wiki/Gary_Miller
Gary Moore	http://en.wikipedia.org/wiki/Gary_Moore
Gary North	http://en.wikipedia.org/wiki/Gary_North_(Christian_Reconstructionist)
Gary Numan	http://en.wikipedia.org/wiki/Gary_Numan
Gary Oldman	http://en.wikipedia.org/wiki/Gary_Oldman
Gary Owens	http://en.wikipedia.org/wiki/Gary_Owens
Gary Peters	http://en.wikipedia.org/wiki/Gary_Peters_(Michigan_politician)
Gary Player	http://en.wikipedia.org/wiki/Gary_Player
Gary Player	http://en.wikipedia.org/wiki/Gary_Player
Gary Ross	http://en.wikipedia.org/wiki/Gary_Ross
Gary Roughead	http://en.wikipedia.org/wiki/Gary_Roughead
Gary S. Becker	http://en.wikipedia.org/wiki/Gary_S._Becker
Gary Sandy	http://en.wikipedia.org/wiki/Gary_Sandy
Gary Sheffield	http://en.wikipedia.org/wiki/Gary_Sheffield
Gary Sinise	http://en.wikipedia.org/wiki/Gary_Sinise
Gary Snyder	http://en.wikipedia.org/wiki/Gary_Snyder
Gary Stevens	http://en.wikipedia.org/wiki/Gary_Stevens
Gary Streeter	http://en.wikipedia.org/wiki/Gary_Streeter
Gary Valentine	http://en.wikipedia.org/wiki/Gary_Valentine
Gary Webb	http://en.wikipedia.org/wiki/Gary_Webb
Gary Wright	http://en.wikipedia.org/wiki/Gary_Wright
Gaspard Bauhin	http://en.wikipedia.org/wiki/Gaspard_Bauhin
Gaston Julia	http://en.wikipedia.org/wiki/Gaston_Julia
Gaston, Duke of Orl�ans	http://en.wikipedia.org/wiki/Gaston%2C_duc_d%27Orl%C3%A9ans
Gates McFadden	http://en.wikipedia.org/wiki/Gates_McFadden
Gavin Arvizo	http://en.wikipedia.org/wiki/Gavin_Arvizo
Gavin Barwell	http://en.wikipedia.org/wiki/Gavin_Barwell
Gavin Bryars	http://en.wikipedia.org/wiki/Gavin_Bryars
Gavin DeGraw	http://en.wikipedia.org/wiki/Gavin_DeGraw
Gavin MacLeod	http://en.wikipedia.org/wiki/Gavin_MacLeod
Gavin Newsom	http://en.wikipedia.org/wiki/Gavin_Newsom
Gavin Rossdale	http://en.wikipedia.org/wiki/Gavin_Rossdale
Gavin Shuker	http://en.wikipedia.org/wiki/Gavin_Shuker
Gavin Williamson	http://en.wikipedia.org/wiki/Gavin_Williamson
Gavriil Derzhavin	http://en.wikipedia.org/wiki/Gavriil_Derzhavin
Gavrilo Princip	http://en.wikipedia.org/wiki/Gavrilo_Princip
Gavyn Davies	http://en.wikipedia.org/wiki/Gavyn_Davies
Gay Talese	http://en.wikipedia.org/wiki/Gay_Talese
Gayatri Spivak	http://en.wikipedia.org/wiki/Gayatri_Spivak
Gayelord Hauser	http://en.wikipedia.org/wiki/Gayelord_Hauser
Gaylord Nelson	http://en.wikipedia.org/wiki/Gaylord_Nelson
Gaylord Perry	http://en.wikipedia.org/wiki/Gaylord_Perry
Gebhard Leberecht von Bl�cher	http://en.wikipedia.org/wiki/Gebhard_Leberecht_von_Bl%C3%Bccher
Gedde Watanabe	http://en.wikipedia.org/wiki/Gedde_Watanabe
Geddy Lee	http://en.wikipedia.org/wiki/Geddy_Lee
G�d�on Tallemant des R�aux	http://en.wikipedia.org/wiki/G%C3%A9d%C3%A9on_Tallemant_des_R%C3%A9aux
Geena Davis	http://en.wikipedia.org/wiki/Geena_Davis
Geezer Butler	http://en.wikipedia.org/wiki/Geezer_Butler
Geir Haarde	http://en.wikipedia.org/wiki/Geir_Haarde
Gelett Burgess	http://en.wikipedia.org/wiki/Gelett_Burgess
Geli Raubal	http://en.wikipedia.org/wiki/Geli_Raubal
Gemma Doyle	http://en.wikipedia.org/wiki/Gemma_Doyle
Gena Rowlands	http://en.wikipedia.org/wiki/Gena_Rowlands
Gene Allison	http://en.wikipedia.org/wiki/Gene_Allison
Gene Anthony Ray	http://en.wikipedia.org/wiki/Gene_Anthony_Ray
Gene Austin	http://en.wikipedia.org/wiki/Gene_Austin
Gene Autry	http://en.wikipedia.org/wiki/Gene_Autry
Gene Barry	http://en.wikipedia.org/wiki/Gene_Barry
Gene Cernan	http://en.wikipedia.org/wiki/Gene_Cernan
Gene Chandler	http://en.wikipedia.org/wiki/Gene_Chandler
Gene Green	http://en.wikipedia.org/wiki/Gene_Green
Gene Hackman	http://en.wikipedia.org/wiki/Gene_Hackman
Gene Kelly	http://en.wikipedia.org/wiki/Gene_Kelly
Gene Krupa	http://en.wikipedia.org/wiki/Gene_Krupa
Gene Lockhart	http://en.wikipedia.org/wiki/Gene_Lockhart
Gene Pitney	http://en.wikipedia.org/wiki/Gene_Pitney
Gene Rayburn	http://en.wikipedia.org/wiki/Gene_Rayburn
Gene Raymond	http://en.wikipedia.org/wiki/Gene_Raymond
Gene Robinson	http://en.wikipedia.org/wiki/Gene_Robinson
Gene Roddenberry	http://en.wikipedia.org/wiki/Gene_Roddenberry
Gene Sarazen	http://en.wikipedia.org/wiki/Gene_Sarazen
Gene Shalit	http://en.wikipedia.org/wiki/Gene_Shalit
Gene Simmons	http://en.wikipedia.org/wiki/Gene_Simmons
Gene Siskel	http://en.wikipedia.org/wiki/Gene_Siskel
Gene Snyder	http://en.wikipedia.org/wiki/Gene_Snyder
Gene Spafford	http://en.wikipedia.org/wiki/Gene_Spafford
Gene Stratton Porter	http://en.wikipedia.org/wiki/Gene_Stratton_Porter
Gene Taylor	http://en.wikipedia.org/wiki/Gene_Taylor_(Mississippi)
Gene Taylor	http://en.wikipedia.org/wiki/Gene_Taylor_(Missouri)
Gene Tierney	http://en.wikipedia.org/wiki/Gene_Tierney
Gene Vincent	http://en.wikipedia.org/wiki/Gene_Vincent
Gene Ween	http://en.wikipedia.org/wiki/Gene_Ween
Gene Wilder	http://en.wikipedia.org/wiki/Gene_Wilder
Gene Wolfe	http://en.wikipedia.org/wiki/Gene_Wolfe
Genesis P-Orridge	http://en.wikipedia.org/wiki/Genesis_P-Orridge
Genevi�ve Bujold	http://en.wikipedia.org/wiki/Genevi%C3%A8ve_Bujold
Genevieve Gorder	http://en.wikipedia.org/wiki/Genevieve_Gorder
Genevieve Taggard	http://en.wikipedia.org/wiki/Genevieve_Taggard
Genghis Khan	http://en.wikipedia.org/wiki/Genghis_Khan
Genie Francis	http://en.wikipedia.org/wiki/Genie_Francis
Gennifer Flowers	http://en.wikipedia.org/wiki/Gennifer_Flowers
Gentile da Fabriano	http://en.wikipedia.org/wiki/Gentile_da_Fabriano
Geoff Barrow	http://en.wikipedia.org/wiki/Geoff_Barrow
Geoff Davis	http://en.wikipedia.org/wiki/Geoff_Davis
Geoff Downes	http://en.wikipedia.org/wiki/Geoff_Downes
Geoff Hoon	http://en.wikipedia.org/wiki/Geoff_Hoon
Geoff Hurst	http://en.wikipedia.org/wiki/Geoff_Hurst
Geoff Rowley	http://en.wikipedia.org/wiki/Geoff_Rowley
Geoff Stults	http://en.wikipedia.org/wiki/Geoff_Stults
Geoffrey Beene	http://en.wikipedia.org/wiki/Geoffrey_Beene
Geoffrey Chaucer	http://en.wikipedia.org/wiki/Geoffrey_Chaucer
Geoffrey Clifton-Brown	http://en.wikipedia.org/wiki/Geoffrey_Clifton-Brown_(born_1953)
Geoffrey Cox	http://en.wikipedia.org/wiki/Geoffrey_Cox
Geoffrey Hartman	http://en.wikipedia.org/wiki/Geoffrey_Hartman
Geoffrey Household	http://en.wikipedia.org/wiki/Geoffrey_Household
Geoffrey Lewis	http://en.wikipedia.org/wiki/Geoffrey_Lewis_(actor)
Geoffrey of Monmouth	http://en.wikipedia.org/wiki/Geoffrey_of_Monmouth
Geoffrey Robinson	http://en.wikipedia.org/wiki/Geoffrey_Robinson
Geoffrey Rowland	http://en.wikipedia.org/wiki/Geoffrey_Rowland
Geoffrey Rush	http://en.wikipedia.org/wiki/Geoffrey_Rush
Geoffrey Wilkinson	http://en.wikipedia.org/wiki/Geoffrey_Wilkinson
Georg Agricola	http://en.wikipedia.org/wiki/Georg_Agricola
Georg B�chner	http://en.wikipedia.org/wiki/Georg_B%C3%Bcchner
Georg Cantor	http://en.wikipedia.org/wiki/Georg_Cantor
Georg Heym	http://en.wikipedia.org/wiki/Georg_Heym
Georg Kaiser	http://en.wikipedia.org/wiki/Georg_Kaiser
Georg Michaelis	http://en.wikipedia.org/wiki/Georg_Michaelis
Georg Philipp Telemann	http://en.wikipedia.org/wiki/Georg_Philipp_Telemann
Georg Rudolf Weckherlin	http://en.wikipedia.org/wiki/Georg_Rudolf_Weckherlin
Georg Simmel	http://en.wikipedia.org/wiki/Georg_Simmel
Georg Simon Ohm	http://en.wikipedia.org/wiki/Georg_Simon_Ohm
Georg Solti	http://en.wikipedia.org/wiki/Georg_Solti
Georg von Hertling	http://en.wikipedia.org/wiki/Georg_von_Hertling
Georg Wilhelm Friedrich Hegel	http://en.wikipedia.org/wiki/Georg_Wilhelm_Friedrich_Hegel
Georg Wittig	http://en.wikipedia.org/wiki/Georg_Wittig
George A. Olah	http://en.wikipedia.org/wiki/George_A._Olah
George A. Parks	http://en.wikipedia.org/wiki/George_A._Parks
George A. Schaefer Jr. 	http://en.wikipedia.org/wiki/George_Schaefer_%28finance%29
George Abbott	http://en.wikipedia.org/wiki/George_Abbott
George Abela	http://en.wikipedia.org/wiki/George_Abela
George Ade	http://en.wikipedia.org/wiki/George_Ade
George Ade	http://en.wikipedia.org/wiki/George_Ade
George Aiken	http://en.wikipedia.org/wiki/George_Aiken
George Akers	http://en.wikipedia.org/wiki/George_Akers
George Akerson	http://en.wikipedia.org/wiki/George_Akerson
George Allen	http://en.wikipedia.org/wiki/George_Allen_(U.S._politician)
George Amy	http://en.wikipedia.org/wiki/George_Amy
George Antheil	http://en.wikipedia.org/wiki/George_Antheil
George Argyros	http://en.wikipedia.org/wiki/George_Argyros
George Arliss	http://en.wikipedia.org/wiki/George_Arliss
George Armstrong Custer	http://en.wikipedia.org/wiki/George_Armstrong_Custer
George B. McClellan	http://en.wikipedia.org/wiki/George_B._McClellan
George B. McClellan, Jr.	http://en.wikipedia.org/wiki/George_B._McClellan%2C_Jr.
George Balanchine	http://en.wikipedia.org/wiki/George_Balanchine
George Bancroft	http://en.wikipedia.org/wiki/George_Bancroft
George Bancroft	http://en.wikipedia.org/wiki/George_Bancroft
George Barker	http://en.wikipedia.org/wiki/George_Barker_(poet)
George Barr McCutcheon	http://en.wikipedia.org/wiki/George_Barr_McCutcheon
George Benson	http://en.wikipedia.org/wiki/George_Benson
George Benson	http://en.wikipedia.org/wiki/George_Benson
George Berkeley	http://en.wikipedia.org/wiki/George_Berkeley
George Bernard Shaw	http://en.wikipedia.org/wiki/George_Bernard_Shaw
George Best	http://en.wikipedia.org/wiki/George_Best
George Biddell Airy	http://en.wikipedia.org/wiki/George_Biddell_Airy
George Blanda	http://en.wikipedia.org/wiki/George_Blanda
George Boole	http://en.wikipedia.org/wiki/George_Boole
George Bowering	http://en.wikipedia.org/wiki/George_Bowering
George Bradshaw	http://en.wikipedia.org/wiki/George_Bradshaw
George Brent	http://en.wikipedia.org/wiki/George_Brent
George Brett	http://en.wikipedia.org/wiki/George_Brett_(baseball)
George Buchanan	http://en.wikipedia.org/wiki/George_Buchanan
George Burns	http://en.wikipedia.org/wiki/George_Burns
George Busbee	http://en.wikipedia.org/wiki/George_Busbee
George Bush	http://en.wikipedia.org/wiki/George_W._Bush
George Busk	http://en.wikipedia.org/wiki/George_Busk
George C. Marshall	http://en.wikipedia.org/wiki/George_C._Marshall
George C. Scott	http://en.wikipedia.org/wiki/George_C._Scott
George C. Wortley	http://en.wikipedia.org/wiki/George_C._Wortley
George Canning	http://en.wikipedia.org/wiki/George_Canning
George Carlin	http://en.wikipedia.org/wiki/George_Carlin
George Cassander	http://en.wikipedia.org/wiki/George_Cassander
George Catlin	http://en.wikipedia.org/wiki/George_Catlin
George Chakiris	http://en.wikipedia.org/wiki/George_Chakiris
George Clinton	http://en.wikipedia.org/wiki/George_Clinton_(musician)
George Clinton	http://en.wikipedia.org/wiki/George_Clinton_(vice_president)
George Clooney	http://en.wikipedia.org/wiki/George_Clooney
George Combe	http://en.wikipedia.org/wiki/George_Combe
George Coulouris	http://en.wikipedia.org/wiki/George_Coulouris
George Creel	http://en.wikipedia.org/wiki/George_Creel
George Cruikshank	http://en.wikipedia.org/wiki/George_Cruikshank
George Crumb	http://en.wikipedia.org/wiki/George_Crumb
George Cukor	http://en.wikipedia.org/wiki/George_Cukor
George Darden	http://en.wikipedia.org/wiki/George_Darden
George Darley	http://en.wikipedia.org/wiki/George_Darley
George David	http://en.wikipedia.org/wiki/George_David
George de Hevesy	http://en.wikipedia.org/wiki/George_de_Hevesy
George Deukmejian	http://en.wikipedia.org/wiki/George_Deukmejian
George Dewey	http://en.wikipedia.org/wiki/George_Dewey
George Douglas	http://en.wikipedia.org/wiki/George_Douglas_Brown
George Douglas Howard Cole	http://en.wikipedia.org/wiki/George_Douglas_Howard_Cole
George du Maurier	http://en.wikipedia.org/wiki/George_du_Maurier
George Duke	http://en.wikipedia.org/wiki/George_Duke
George Dzundza	http://en.wikipedia.org/wiki/George_Dzundza
George E. Brown, Jr.	http://en.wikipedia.org/wiki/George_E._Brown%2C_Jr.
George E. MacKinnon	http://en.wikipedia.org/wiki/George_E._MacKinnon
George E. Marshall	http://en.wikipedia.org/wiki/George_Marshall_%28director%29
George E. Reedy	http://en.wikipedia.org/wiki/George_E._Reedy
George Eads	http://en.wikipedia.org/wiki/George_Eads
George Eastman	http://en.wikipedia.org/wiki/George_Eastman
George Edmund Street	http://en.wikipedia.org/wiki/George_Edmund_Street
George Eliot	http://en.wikipedia.org/wiki/George_Eliot
George Ellery Hale	http://en.wikipedia.org/wiki/George_Ellery_Hale
George Etherege	http://en.wikipedia.org/wiki/George_Etherege
George Eustice	http://en.wikipedia.org/wiki/George_Eustice
George Evans	http://en.wikipedia.org/wiki/George_Evans_%28comics%29
George F. Kennan	http://en.wikipedia.org/wiki/George_F._Kennan
George Farquhar	http://en.wikipedia.org/wiki/George_Farquhar
George Foreman	http://en.wikipedia.org/wiki/George_Foreman
George Frederick Baer	http://en.wikipedia.org/wiki/George_Frederick_Baer
George Freeman	http://en.wikipedia.org/wiki/George_Freeman_(politician)
George Frideric Handel	http://en.wikipedia.org/wiki/George_Frideric_Handel
George Gabriel Stokes	http://en.wikipedia.org/wiki/George_Gabriel_Stokes
George Galloway	http://en.wikipedia.org/wiki/George_Galloway
George Gallup	http://en.wikipedia.org/wiki/George_Gallup
George Gamow	http://en.wikipedia.org/wiki/George_Gamow
George Gaynes	http://en.wikipedia.org/wiki/George_Gaynes
George Gershwin	http://en.wikipedia.org/wiki/George_Gershwin
George Gilder	http://en.wikipedia.org/wiki/George_Gilder
George Gissing	http://en.wikipedia.org/wiki/George_Gissing
George Gobel	http://en.wikipedia.org/wiki/George_Gobel
George Goethals	http://en.wikipedia.org/wiki/George_Goethals
George Gordon Meade	http://en.wikipedia.org/wiki/George_Gordon_Meade
George Grenville	http://en.wikipedia.org/wiki/George_Grenville
George Grossmith	http://en.wikipedia.org/wiki/George_Grossmith
George Grosz	http://en.wikipedia.org/wiki/George_Grosz
George H. Fallon	http://en.wikipedia.org/wiki/George_H._Fallon
George H.W. Bush	http://en.wikipedia.org/wiki/George_H.W._Bush
George Halas	http://en.wikipedia.org/wiki/George_Halas
George Hamilton	http://en.wikipedia.org/wiki/George_Hamilton_(actor)
George Harrison	http://en.wikipedia.org/wiki/George_Harrison
George Hennard	http://en.wikipedia.org/wiki/George_Hennard
George Henry Boker	http://en.wikipedia.org/wiki/George_Henry_Boker
George Henry Lewes	http://en.wikipedia.org/wiki/George_Henry_Lewes
George Henry Thomas	http://en.wikipedia.org/wiki/George_Henry_Thomas
George Herbert	http://en.wikipedia.org/wiki/George_Herbert
George Herbert Mead	http://en.wikipedia.org/wiki/George_Herbert_Mead
George Herbert Walker III	http://en.wikipedia.org/wiki/George_Herbert_Walker_III
George Hickes	http://en.wikipedia.org/wiki/George_Hickes
George Hollingbery	http://en.wikipedia.org/wiki/George_Hollingbery
George Howarth	http://en.wikipedia.org/wiki/George_Howarth
George Inness	http://en.wikipedia.org/wiki/George_Inness
George J. Mitchell	http://en.wikipedia.org/wiki/George_J._Mitchell
George J. Mitchell	http://en.wikipedia.org/wiki/George_J._Mitchell
George J. Stigler	http://en.wikipedia.org/wiki/George_J._Stigler
George James Symons	http://en.wikipedia.org/wiki/George_James_Symons
George Jean Nathan	http://en.wikipedia.org/wiki/George_Jean_Nathan
George Jones	http://en.wikipedia.org/wiki/George_Jones
George Jung	http://en.wikipedia.org/wiki/George_Jung
George Kelly	http://en.wikipedia.org/wiki/George_Kelly_(playwright)
George Kennedy	http://en.wikipedia.org/wiki/George_Kennedy
George L. Aiken	http://en.wikipedia.org/wiki/George_Aiken_%28playwright%29
George Lazenby	http://en.wikipedia.org/wiki/George_Lazenby
George LeMieux	http://en.wikipedia.org/wiki/George_LeMieux
George Lindsey	http://en.wikipedia.org/wiki/George_Lindsey
George Lopez	http://en.wikipedia.org/wiki/George_Lopez
George Lucas	http://en.wikipedia.org/wiki/George_Lucas
George M. Cohan	http://en.wikipedia.org/wiki/George_M._Cohan
George M. Dallas	http://en.wikipedia.org/wiki/George_M._Dallas
George M. O'Brien	http://en.wikipedia.org/wiki/George_M._O%27Brien
George MacDonald	http://en.wikipedia.org/wiki/George_MacDonald
George Maciunas	http://en.wikipedia.org/wiki/George_Maciunas
George Mackay Brown	http://en.wikipedia.org/wiki/George_Mackay_Brown
George Macready	http://en.wikipedia.org/wiki/George_Macready
George Maharis	http://en.wikipedia.org/wiki/George_Maharis
George Mallory	http://en.wikipedia.org/wiki/George_Mallory
George Martin	http://en.wikipedia.org/wiki/George_Martin
George Mason	http://en.wikipedia.org/wiki/George_Mason
George Maxwell Richards	http://en.wikipedia.org/wiki/George_Maxwell_Richards
George McDuffie	http://en.wikipedia.org/wiki/George_McDuffie
George McGovern	http://en.wikipedia.org/wiki/George_McGovern
George Meany	http://en.wikipedia.org/wiki/George_Meany
George Meredith	http://en.wikipedia.org/wiki/George_Meredith
George Michael	http://en.wikipedia.org/wiki/George_Michael
George Mikan	http://en.wikipedia.org/wiki/George_Mikan
George Miller	http://en.wikipedia.org/wiki/George_Miller_(California_politician)
George Miller	http://en.wikipedia.org/wiki/George_Miller,_Jr.
George Montgomery	http://en.wikipedia.org/wiki/George_Montgomery
George Morfogen	http://en.wikipedia.org/wiki/George_Morfogen
George Moscone	http://en.wikipedia.org/wiki/George_Moscone
George Moses Horton	http://en.wikipedia.org/wiki/George_Moses_Horton
George Mudie	http://en.wikipedia.org/wiki/George_Mudie
George Murphy	http://en.wikipedia.org/wiki/George_Murphy
George Nader	http://en.wikipedia.org/wiki/George_Nader
George Nethercutt	http://en.wikipedia.org/wiki/George_Nethercutt
George Oppen	http://en.wikipedia.org/wiki/George_Oppen
George Orwell	http://en.wikipedia.org/wiki/George_Orwell
George Osborne	http://en.wikipedia.org/wiki/George_Osborne
George Packer	http://en.wikipedia.org/wiki/George_Packer
George Paget Thomson	http://en.wikipedia.org/wiki/George_Paget_Thomson
George Pake	http://en.wikipedia.org/wiki/George_Pake
George Pal	http://en.wikipedia.org/wiki/George_Pal
George Papandreou	http://en.wikipedia.org/wiki/George_Papandreou_(junior)
George Pataki	http://en.wikipedia.org/wiki/George_Pataki
George Pataki	http://en.wikipedia.org/wiki/George_Pataki
George Payne Rainsford James	http://en.wikipedia.org/wiki/George_Payne_Rainsford_James
George Peabody	http://en.wikipedia.org/wiki/George_Peabody
George Peacock	http://en.wikipedia.org/wiki/George_Peacock
George Peele	http://en.wikipedia.org/wiki/George_Peele
George Peppard	http://en.wikipedia.org/wiki/George_Peppard
George Plimpton	http://en.wikipedia.org/wiki/George_Plimpton
George Porter	http://en.wikipedia.org/wiki/George_Porter
George Pullman	http://en.wikipedia.org/wiki/George_Pullman
George Puttenham	http://en.wikipedia.org/wiki/George_Puttenham
George R. R. Martin	http://en.wikipedia.org/wiki/George_R._R._Martin
George Radanovich	http://en.wikipedia.org/wiki/George_Radanovich
George Raft	http://en.wikipedia.org/wiki/George_Raft
George Reeves	http://en.wikipedia.org/wiki/George_Reeves
George Ripley	http://en.wikipedia.org/wiki/George_Ripley_%28transcendentalist%29
George Rockwell	http://en.wikipedia.org/wiki/George_Rockwell
George Rogers Clark	http://en.wikipedia.org/wiki/George_Rogers_Clark
George Romero	http://en.wikipedia.org/wiki/George_Romero
George Roy Hill	http://en.wikipedia.org/wiki/George_Roy_Hill
George Ryan	http://en.wikipedia.org/wiki/George_Ryan
George S. Kaufman	http://en.wikipedia.org/wiki/George_S._Kaufman
George S. Patton	http://en.wikipedia.org/wiki/George_S._Patton
George Saintsbury	http://en.wikipedia.org/wiki/George_Saintsbury
George Sand	http://en.wikipedia.org/wiki/George_Sand
George Sanders	http://en.wikipedia.org/wiki/George_Sanders
George Santayana	http://en.wikipedia.org/wiki/George_Santayana
George Sarton	http://en.wikipedia.org/wiki/George_Sarton
George Segal	http://en.wikipedia.org/wiki/George_Segal
George Shultz	http://en.wikipedia.org/wiki/George_Shultz
George Sidney	http://en.wikipedia.org/wiki/George_Sidney
George Sisler	http://en.wikipedia.org/wiki/George_Sisler
George Smathers	http://en.wikipedia.org/wiki/George_Smathers
George Soros	http://en.wikipedia.org/wiki/George_Soros
George Steinbrenner	http://en.wikipedia.org/wiki/George_Steinbrenner
George Steiner	http://en.wikipedia.org/wiki/George_Steiner
George Stephanopoulos	http://en.wikipedia.org/wiki/George_Stephanopoulos
George Stephenson	http://en.wikipedia.org/wiki/George_Stephenson
George Stevens	http://en.wikipedia.org/wiki/George_Stevens
George Stoneman	http://en.wikipedia.org/wiki/George_Stoneman
George Strait	http://en.wikipedia.org/wiki/George_Strait
George Stults	http://en.wikipedia.org/wiki/George_Stults
George Takei	http://en.wikipedia.org/wiki/George_Takei
George Tenet	http://en.wikipedia.org/wiki/George_Tenet
George Thorogood	http://en.wikipedia.org/wiki/George_Thorogood
George Ticknor	http://en.wikipedia.org/wiki/George_Ticknor
George Ticknor Curtis	http://en.wikipedia.org/wiki/George_Ticknor_Curtis
George Uhlenbeck	http://en.wikipedia.org/wiki/George_Uhlenbeck
George Vancouver	http://en.wikipedia.org/wiki/George_Vancouver
George Vasiliou	http://en.wikipedia.org/wiki/George_Vasiliou
George Voinovich	http://en.wikipedia.org/wiki/George_Voinovich
George W. Bush	http://en.wikipedia.org/wiki/George_W._Bush
George W. Cable	http://en.wikipedia.org/wiki/George_W._Cable
George W. Crockett, Jr.	http://en.wikipedia.org/wiki/George_W._Crockett%2C_Jr.
George W. Gekas	http://en.wikipedia.org/wiki/George_W._Gekas
George W. Romney	http://en.wikipedia.org/wiki/George_W._Romney
George Wackenhut	http://en.wikipedia.org/wiki/George_Wackenhut
George Wald	http://en.wikipedia.org/wiki/George_Wald
George Wallace	http://en.wikipedia.org/wiki/George_Wallace
George Washington	http://en.wikipedia.org/wiki/George_Washington
George Washington Carver	http://en.wikipedia.org/wiki/George_Washington_Carver
George Washington Owen	http://en.wikipedia.org/wiki/George_Washington_Owen
George Weah	http://en.wikipedia.org/wiki/George_Weah
George Wendt	http://en.wikipedia.org/wiki/George_Wendt
George Westinghouse	http://en.wikipedia.org/wiki/George_Westinghouse
George White	http://en.wikipedia.org/wiki/George_White_(Ohio_politician)
George Whitefield	http://en.wikipedia.org/wiki/George_Whitefield
George Will	http://en.wikipedia.org/wiki/George_Will
George Wishart	http://en.wikipedia.org/wiki/George_Wishart
George Young	http://en.wikipedia.org/wiki/Sir_George_Young,_6th_Baronet
George Zoley	http://en.wikipedia.org/wiki/George_Zoley
Georges Auric	http://en.wikipedia.org/wiki/Georges_Auric
Georges Bataille	http://en.wikipedia.org/wiki/Georges_Bataille
Georges Bernanos	http://en.wikipedia.org/wiki/Georges_Bernanos
Georges Bizet	http://en.wikipedia.org/wiki/Georges_Bizet
Georges Braque	http://en.wikipedia.org/wiki/Georges_Braque
Georges Charpak	http://en.wikipedia.org/wiki/Georges_Charpak
Georges Clemenceau	http://en.wikipedia.org/wiki/Georges_Clemenceau
Georges Cuvier	http://en.wikipedia.org/wiki/Georges_Cuvier
Georges d'Amboise	http://en.wikipedia.org/wiki/Georges_d%27Amboise
Georges Delerue	http://en.wikipedia.org/wiki/Georges_Delerue
Georges Duhamel	http://en.wikipedia.org/wiki/Georges_Duhamel
Georges Jacques Danton	http://en.wikipedia.org/wiki/Georges_Jacques_Danton
Georges Perec	http://en.wikipedia.org/wiki/Georges_Perec
Georges Pire	http://en.wikipedia.org/wiki/Georges_Pire
Georges Pompidou	http://en.wikipedia.org/wiki/Georges_Pompidou
Georges Rouault	http://en.wikipedia.org/wiki/Georges_Rouault
Georges Seurat	http://en.wikipedia.org/wiki/Georges_Seurat
Georges Simenon	http://en.wikipedia.org/wiki/Georges_Simenon
Georges-Louis Leclerc, Comte de Buffon	http://en.wikipedia.org/wiki/Georges-Louis_Leclerc%2C_Comte_de_Buffon
Georgi Djulgerov	http://en.wikipedia.org/wiki/Georgi_Djulgerov
Georgi Markov	http://en.wikipedia.org/wiki/Georgi_Markov
Georgi Parvanov	http://en.wikipedia.org/wiki/Georgi_Parvanov
Georgi Zhukov	http://en.wikipedia.org/wiki/Georgi_Zhukov
Georgia Brown	http://en.wikipedia.org/wiki/Georgia_Brown_(English_singer)
Georgia O'Keeffe	http://en.wikipedia.org/wiki/Georgia_O%27Keeffe
Georgie Fame	http://en.wikipedia.org/wiki/Georgie_Fame
Georgius Macropedius	http://en.wikipedia.org/wiki/Georgius_Macropedius
Geraint Davies	http://en.wikipedia.org/wiki/Geraint_Davies_%28Labour_politician%29
Gerald A. Soffen	http://en.wikipedia.org/wiki/Gerald_Soffen
Gerald B.H. Solomon	http://en.wikipedia.org/wiki/Gerald_B.H._Solomon
Gerald Casale	http://en.wikipedia.org/wiki/Gerald_Casale
Gerald D. Kleczka	http://en.wikipedia.org/wiki/Gerald_D._Kleczka
Gerald Durrell	http://en.wikipedia.org/wiki/Gerald_Durrell
Gerald Ford	http://en.wikipedia.org/wiki/Gerald_Ford
Gerald Gardner	http://en.wikipedia.org/wiki/Gerald_Gardner
Gerald Howarth	http://en.wikipedia.org/wiki/Gerald_Howarth
Gerald Kaufman	http://en.wikipedia.org/wiki/Gerald_Kaufman
Gerald L. Baliles	http://en.wikipedia.org/wiki/Gerald_L._Baliles
Gerald McRaney	http://en.wikipedia.org/wiki/Gerald_McRaney
Geraldine Brooks	http://en.wikipedia.org/wiki/Geraldine_Brooks_(writer)
Geraldine Chaplin	http://en.wikipedia.org/wiki/Geraldine_Chaplin
Geraldine Ferraro	http://en.wikipedia.org/wiki/Geraldine_Ferraro
Geraldine Fitzgerald	http://en.wikipedia.org/wiki/Geraldine_Fitzgerald
Geraldine Laybourne	http://en.wikipedia.org/wiki/Geraldine_Laybourne
Geraldine Page	http://en.wikipedia.org/wiki/Geraldine_Page
Geraldo Rivera	http://en.wikipedia.org/wiki/Geraldo_Rivera
Gerard Arpey	http://en.wikipedia.org/wiki/Gerard_Arpey
Gerard Butler	http://en.wikipedia.org/wiki/Gerard_Butler
Gerard David	http://en.wikipedia.org/wiki/Gerard_David
G�rard de Nerval	http://en.wikipedia.org/wiki/G%C3%A9rard_de_Nerval
Gerard Depardieu	http://en.wikipedia.org/wiki/Gerard_Depardieu
G�rard Latortue	http://en.wikipedia.org/wiki/G%C3%A9rard_Latortue
Gerard Manley Hopkins	http://en.wikipedia.org/wiki/Gerard_Manley_Hopkins
Gerard Mercator	http://en.wikipedia.org/wiki/Gerard_Mercator
G�rard Paul Deshayes	http://en.wikipedia.org/wiki/G%C3%A9rard_Paul_Deshayes
Gerard Terborch	http://en.wikipedia.org/wiki/Gerard_Terborch
Gerard Way	http://en.wikipedia.org/wiki/Gerard_Way
Gerardus 't Hooft	http://en.wikipedia.org/wiki/Gerardus_%27t_Hooft
Gerbrand van den Eeckhout	http://en.wikipedia.org/wiki/Gerbrand_van_den_Eeckhout
Gerd Binnig	http://en.wikipedia.org/wiki/Gerd_Binnig
Gerd Muller	http://en.wikipedia.org/wiki/Gerd_Muller
Gerd von Rundstedt	http://en.wikipedia.org/wiki/Gerd_von_Rundstedt
Gerhard Herzberg	http://en.wikipedia.org/wiki/Gerhard_Herzberg
Gerhard Schroeder	http://en.wikipedia.org/wiki/Gerhard_Schroeder
Gerhart Hauptmann	http://en.wikipedia.org/wiki/Gerhart_Hauptmann
Geri Halliwell	http://en.wikipedia.org/wiki/Geri_Halliwell
Germaine Greer	http://en.wikipedia.org/wiki/Germaine_Greer
Germaine Tailleferre	http://en.wikipedia.org/wiki/Germaine_Tailleferre
Germanicus Caesar	http://en.wikipedia.org/wiki/Germanicus_Caesar
Gerrit Smith	http://en.wikipedia.org/wiki/Gerrit_Smith
Gerrit van Honthorst	http://en.wikipedia.org/wiki/Gerrit_van_Honthorst
Gerry Adams	http://en.wikipedia.org/wiki/Gerry_Adams
Gerry Beckley	http://en.wikipedia.org/wiki/Gerry_Beckley
Gerry Connolly	http://en.wikipedia.org/wiki/Gerry_Connolly
Gerry Cooney	http://en.wikipedia.org/wiki/Gerry_Cooney
Gerry E. Studds	http://en.wikipedia.org/wiki/Gerry_E._Studds
Gerry McCambridge	http://en.wikipedia.org/wiki/Gerry_McCambridge
Gerry Mulligan	http://en.wikipedia.org/wiki/Gerry_Mulligan
Gerry Sikorski	http://en.wikipedia.org/wiki/Gerry_Sikorski
Gerry Studds	http://en.wikipedia.org/wiki/Gerry_Studds
Gerry Sutcliffe	http://en.wikipedia.org/wiki/Gerry_Sutcliffe
Gertrude Himmelfarb	http://en.wikipedia.org/wiki/Gertrude_Himmelfarb
Gertrude Lawrence	http://en.wikipedia.org/wiki/Gertrude_Lawrence
Gertrude Stein	http://en.wikipedia.org/wiki/Gertrude_Stein
Gertrude Vanderbilt Whitney	http://en.wikipedia.org/wiki/Gertrude_Vanderbilt_Whitney
Get�lio Vargas	http://en.wikipedia.org/wiki/Get%C3%BAlio_Vargas
Ghazi al-Yawar	http://en.wikipedia.org/wiki/Ghazi_al-Yawar
Ghostface Killah	http://en.wikipedia.org/wiki/Ghostface_Killah
Gia Carangi	http://en.wikipedia.org/wiki/Gia_Carangi
Giacomo Agostini	http://en.wikipedia.org/wiki/Giacomo_Agostini
Giacomo Casanova	http://en.wikipedia.org/wiki/Giacomo_Casanova
Giacomo Leopardi	http://en.wikipedia.org/wiki/Giacomo_Leopardi
Giacomo Meyerbeer	http://en.wikipedia.org/wiki/Giacomo_Meyerbeer
Giacomo Puccini	http://en.wikipedia.org/wiki/Giacomo_Puccini
Giambattista Bodoni	http://en.wikipedia.org/wiki/Giambattista_Bodoni
Giambattista della Porta	http://en.wikipedia.org/wiki/Giambattista_della_Porta
Giambattista Piranesi	http://en.wikipedia.org/wiki/Giambattista_Piranesi
Gian Francesco Malipiero	http://en.wikipedia.org/wiki/Gian_Francesco_Malipiero
Gian Lorenzo Bernini	http://en.wikipedia.org/wiki/Gian_Lorenzo_Bernini
Giancarlo Esposito	http://en.wikipedia.org/wiki/Giancarlo_Esposito
Gian-Carlo Menotti	http://en.wikipedia.org/wiki/Gian-Carlo_Menotti
Gianfranco Zola	http://en.wikipedia.org/wiki/Gianfranco_Zola
Giangiorgio Trissino	http://en.wikipedia.org/wiki/Giangiorgio_Trissino
Gianni Agnelli	http://en.wikipedia.org/wiki/Gianni_Agnelli
Gianni Vattimo	http://en.wikipedia.org/wiki/Gianni_Vattimo
Gianni Versace	http://en.wikipedia.org/wiki/Gianni_Versace
Gideon Mantell	http://en.wikipedia.org/wiki/Gideon_Mantell
Gig Young	http://en.wikipedia.org/wiki/Gig_Young
Gijs de Vries	http://en.wikipedia.org/wiki/Gijs_de_Vries
Gil Amelio	http://en.wikipedia.org/wiki/Gil_Amelio
Gil Bellows	http://en.wikipedia.org/wiki/Gil_Bellows
Gil Evans	http://en.wikipedia.org/wiki/Gil_Evans
Gil Gerard	http://en.wikipedia.org/wiki/Gil_Gerard
Gil Gutknecht	http://en.wikipedia.org/wiki/Gil_Gutknecht
Gil Hodges	http://en.wikipedia.org/wiki/Gil_Hodges
Gil Kerlikowske	http://en.wikipedia.org/wiki/Gil_Kerlikowske
Gilbert Amy	http://en.wikipedia.org/wiki/Gilbert_Amy
Gilbert Burnet	http://en.wikipedia.org/wiki/Gilbert_Burnet
Gilbert de la Porr�e	http://en.wikipedia.org/wiki/Gilbert_de_la_Porr%C3%A9e
Gilbert Gottfried	http://en.wikipedia.org/wiki/Gilbert_Gottfried
Gilbert Hernandez	http://en.wikipedia.org/wiki/Gilbert_Gottfried
Gilbert Houngbo	http://en.wikipedia.org/wiki/Gilbert_Houngbo
Gilbert M. Anderson	http://en.wikipedia.org/wiki/Gilbert_M._Anderson
Gilbert Roland	http://en.wikipedia.org/wiki/Gilbert_Roland
Gilbert Sheldon	http://en.wikipedia.org/wiki/Gilbert_Sheldon
Gilbert Stuart	http://en.wikipedia.org/wiki/Gilbert_Stuart
Gilbert White	http://en.wikipedia.org/wiki/Gilbert_White
Gilda Radner	http://en.wikipedia.org/wiki/Gilda_Radner
Gilles de Rais	http://en.wikipedia.org/wiki/Gilles_de_Rais
Gilles Personne de Roberval	http://en.wikipedia.org/wiki/Gilles_Personne_de_Roberval
Gillian Anderson	http://en.wikipedia.org/wiki/Gillian_Anderson
Gillian Armstrong	http://en.wikipedia.org/wiki/Gillian_Armstrong
Gina Albert	http://en.wikipedia.org/wiki/Gina_Albert
Gina Gershon	http://en.wikipedia.org/wiki/Gina_Gershon
Gina Lollobrigida	http://en.wikipedia.org/wiki/Gina_Lollobrigida
Gina Philips	http://en.wikipedia.org/wiki/Gina_Philips
Gina Schock	http://en.wikipedia.org/wiki/Gina_Schock
Gina Torres	http://en.wikipedia.org/wiki/Gina_Torres
Ginger Baker	http://en.wikipedia.org/wiki/Ginger_Baker
Ginger Rogers	http://en.wikipedia.org/wiki/Ginger_Rogers
Ginnifer Goodwin	http://en.wikipedia.org/wiki/Ginnifer_Goodwin
Ginny Brown-Waite	http://en.wikipedia.org/wiki/Ginny_Brown-Waite
Gioacchino Rossini	http://en.wikipedia.org/wiki/Gioacchino_Rossini
Gioconda Belli	http://en.wikipedia.org/wiki/Gioconda_Belli
Giordano Bruno	http://en.wikipedia.org/wiki/Giordano_Bruno
Giorgio Armani	http://en.wikipedia.org/wiki/Giorgio_Armani
Giorgio de Chirico	http://en.wikipedia.org/wiki/Giorgio_de_Chirico
Giorgio Moroder	http://en.wikipedia.org/wiki/Giorgio_Moroder
Giorgio Napolitano	http://en.wikipedia.org/wiki/Giorgio_Napolitano
Giorgio Vasari	http://en.wikipedia.org/wiki/Giorgio_Vasari
Giorgos Seferis	http://en.wikipedia.org/wiki/Giorgos_Seferis
Giosu� Carducci	http://en.wikipedia.org/wiki/Giosu%C3%A8_Carducci
Giotto di Bondone	http://en.wikipedia.org/wiki/Giotto_di_Bondone
Giovanni Alfonso Borelli	http://en.wikipedia.org/wiki/Giovanni_Alfonso_Borelli
Giovanni Battista Amici	http://en.wikipedia.org/wiki/Giovanni_Battista_Amici
Giovanni Battista Casti	http://en.wikipedia.org/wiki/Giovanni_Battista_Casti
Giovanni Battista Pergolesi	http://en.wikipedia.org/wiki/Giovanni_Battista_Pergolesi
Giovanni Battista Tiepolo	http://en.wikipedia.org/wiki/Giovanni_Battista_Tiepolo
Giovanni Bellini	http://en.wikipedia.org/wiki/Giovanni_Bellini
Giovanni Benedetto Castiglione	http://en.wikipedia.org/wiki/Giovanni_Benedetto_Castiglione
Giovanni Boccaccio	http://en.wikipedia.org/wiki/Giovanni_Boccaccio
Giovanni Bottesini	http://en.wikipedia.org/wiki/Giovanni_Bottesini
Giovanni da Verrazano	http://en.wikipedia.org/wiki/Giovanni_da_Verrazano
Giovanni Della Casa	http://en.wikipedia.org/wiki/Giovanni_Della_Casa
Giovanni Domenico Cassini	http://en.wikipedia.org/wiki/Giovanni_Domenico_Cassini
Giovanni Gabrieli	http://en.wikipedia.org/wiki/Giovanni_Gabrieli
Giovanni Paisiello	http://en.wikipedia.org/wiki/Giovanni_Paisiello
Giovanni Pico della Mirandola	http://en.wikipedia.org/wiki/Giovanni_Pico_della_Mirandola
Giovanni Pierluigi da Palestrina	http://en.wikipedia.org/wiki/Giovanni_Pierluigi_da_Palestrina
Giovanni Pisano	http://en.wikipedia.org/wiki/Giovanni_Pisano
Giovanni Ribisi	http://en.wikipedia.org/wiki/Giovanni_Ribisi
Giovanni Virginio Schiaparelli	http://en.wikipedia.org/wiki/Giovanni_Virginio_Schiaparelli
Girija Prasad Koirala	http://en.wikipedia.org/wiki/Girija_Prasad_Koirala
Girma Wolde-Giorgis	http://en.wikipedia.org/wiki/Girma_Wolde-Giorgis
Girolamo Cardano	http://en.wikipedia.org/wiki/Girolamo_Cardano
Girolamo Fabrici	http://en.wikipedia.org/wiki/Girolamo_Fabrici
Girolamo Frescobaldi	http://en.wikipedia.org/wiki/Girolamo_Frescobaldi
Girolamo Muziano	http://en.wikipedia.org/wiki/Girolamo_Muziano
Girolamo Savonarola	http://en.wikipedia.org/wiki/Girolamo_Savonarola
Gisela Stuart	http://en.wikipedia.org/wiki/Gisela_Stuart
Gisele Bundchen	http://en.wikipedia.org/wiki/Gisele_Bundchen
Giuliana Sgrena	http://en.wikipedia.org/wiki/Giuliana_Sgrena
Giulio Alberoni	http://en.wikipedia.org/wiki/Giulio_Alberoni
Giulio Andreotti	http://en.wikipedia.org/wiki/Giulio_Andreotti
Giulio Douhet	http://en.wikipedia.org/wiki/Giulio_Douhet
Giulio Natta	http://en.wikipedia.org/wiki/Giulio_Natta
Giulio Romano	http://en.wikipedia.org/wiki/Giulio_Romano
Giuseppe Addobbati	http://en.wikipedia.org/wiki/Giuseppe_Addobbati
Giuseppe Alizeri	http://en.wikipedia.org/wiki/Giuseppe_Alizeri
Giuseppe Arcimboldo	http://en.wikipedia.org/wiki/Giuseppe_Arcimboldo
Giuseppe Garibaldi	http://en.wikipedia.org/wiki/Giuseppe_Garibaldi
Giuseppe Marco Fieschi	http://en.wikipedia.org/wiki/Giuseppe_Marco_Fieschi
Giuseppe Maria Crespi	http://en.wikipedia.org/wiki/Giuseppe_Maria_Crespi
Giuseppe Mazzini	http://en.wikipedia.org/wiki/Giuseppe_Mazzini
Giuseppe Parini	http://en.wikipedia.org/wiki/Giuseppe_Parini
Giuseppe Peano	http://en.wikipedia.org/wiki/Giuseppe_Peano
Giuseppe Sarti	http://en.wikipedia.org/wiki/Giuseppe_Sarti
Giuseppe Tartini	http://en.wikipedia.org/wiki/Giuseppe_Tartini
Giuseppe Tomasi di Lampedusa	http://en.wikipedia.org/wiki/Giuseppe_Tomasi_di_Lampedusa
Giuseppe Verdi	http://en.wikipedia.org/wiki/Giuseppe_Verdi
Giuseppe Zangara	http://en.wikipedia.org/wiki/Giuseppe_Zangara
Gjorge Ivanov	http://en.wikipedia.org/wiki/Gjorge_Ivanov
Gladwyn Jebb	http://en.wikipedia.org/wiki/Gladwyn_Jebb
Gladys Knight	http://en.wikipedia.org/wiki/Gladys_Knight
Glen Campbell	http://en.wikipedia.org/wiki/Glen_Campbell
Glen E. Edgerton	http://en.wikipedia.org/wiki/Glen_E._Edgerton
Glen Matlock	http://en.wikipedia.org/wiki/Glen_Matlock
Glenda Hood	http://en.wikipedia.org/wiki/Glenda_Hood
Glenda Jackson	http://en.wikipedia.org/wiki/Glenda_Jackson
Glenn Beck	http://en.wikipedia.org/wiki/Glenn_Beck
Glenn Close	http://en.wikipedia.org/wiki/Glenn_Close
Glenn Curtiss	http://en.wikipedia.org/wiki/Glenn_Curtiss
Glenn Danzig	http://en.wikipedia.org/wiki/Glenn_Danzig
Glenn English	http://en.wikipedia.org/wiki/Glenn_English
Glenn English	http://en.wikipedia.org/wiki/Glenn_English
Glenn Ford	http://en.wikipedia.org/wiki/Glenn_Ford
Glenn Frey	http://en.wikipedia.org/wiki/Glenn_Frey
Glenn Gould	http://en.wikipedia.org/wiki/Glenn_Gould
Glenn Hoddle	http://en.wikipedia.org/wiki/Glenn_Hoddle
Glenn Hubbard	http://en.wikipedia.org/wiki/Glenn_Hubbard_(economics)
Glenn M. Anderson	http://en.wikipedia.org/wiki/Glenn_M._Anderson
Glenn Miller	http://en.wikipedia.org/wiki/Glenn_Miller
Glenn Nye	http://en.wikipedia.org/wiki/Glenn_Nye
Glenn Quinn	http://en.wikipedia.org/wiki/Glenn_Quinn
Glenn Seaborg	http://en.wikipedia.org/wiki/Glenn_Seaborg
Glenn Thompson	http://en.wikipedia.org/wiki/Glenn_
Glenne Headly	http://en.wikipedia.org/wiki/Glenne_Headly
Glenway Wescott	http://en.wikipedia.org/wiki/Glenway_Wescott
Gloria Allred	http://en.wikipedia.org/wiki/Gloria_Allred
Gloria De Piero	http://en.wikipedia.org/wiki/Gloria_De_Piero
Gloria DeHaven	http://en.wikipedia.org/wiki/Gloria_DeHaven
Gloria Dickson	http://en.wikipedia.org/wiki/Gloria_Dickson
Gloria Estefan	http://en.wikipedia.org/wiki/Gloria_Estefan
Gloria Gaynor	http://en.wikipedia.org/wiki/Gloria_Gaynor
Gloria Grahame	http://en.wikipedia.org/wiki/Gloria_Grahame
Gloria Macapagal-Arroyo	http://en.wikipedia.org/wiki/Gloria_Macapagal-Arroyo
Gloria Macapagal-Arroyo	http://en.wikipedia.org/wiki/Gloria_Macapagal-Arroyo
Gloria Naylor	http://en.wikipedia.org/wiki/Gloria_Naylor
Gloria Reuben	http://en.wikipedia.org/wiki/Gloria_Reuben
Gloria Steinem	http://en.wikipedia.org/wiki/Gloria_Steinem
Gloria Stuart	http://en.wikipedia.org/wiki/Gloria_Stuart
Gloria Swanson	http://en.wikipedia.org/wiki/Gloria_Swanson
Gloria Trevi	http://en.wikipedia.org/wiki/Gloria_Trevi
Gloria Tristani	http://en.wikipedia.org/wiki/Gloria_Tristani
Gloria Vanderbilt	http://en.wikipedia.org/wiki/Gloria_Vanderbilt
Glyn Davies	http://en.wikipedia.org/wiki/Glyn_Davies_(Welsh_politician)
Gnassingbe Eyadema	http://en.wikipedia.org/wiki/Gnassingbe_Eyadema
Godfrey Cambridge	http://en.wikipedia.org/wiki/Godfrey_Cambridge
Godfrey Reggio	http://en.wikipedia.org/wiki/Godfrey_Reggio
Godfried Danneels	http://en.wikipedia.org/wiki/Godfried_Danneels
Gogi Grant	http://en.wikipedia.org/wiki/Gogi_Grant
Goh Chok Tong	http://en.wikipedia.org/wiki/Goh_Chok_Tong
Gold Chains	http://en.wikipedia.org/wiki/Gold_Chains
Golda Meir	http://en.wikipedia.org/wiki/Golda_Meir
Golden Brooks	http://en.wikipedia.org/wiki/Golden_Brooks
Goldie Hawn	http://en.wikipedia.org/wiki/Goldie_Hawn
Goldy McJohn	http://en.wikipedia.org/wiki/Goldy_McJohn
Gong Li	http://en.wikipedia.org/wiki/Gong_Li
Gonzalo de C�spedes y Meneses	http://en.wikipedia.org/wiki/Gonzalo_de_C%C3%A9spedes_y_Meneses
Goodluck Jonathan	http://en.wikipedia.org/wiki/Goodluck_Jonathan
Goodman Ace	http://en.wikipedia.org/wiki/Goodman_Ace
Googie Withers	http://en.wikipedia.org/wiki/Googie_Withers
G�ran Persson	http://en.wikipedia.org/wiki/G%C3%B6ran_Persson
Goran Visnjic	http://en.wikipedia.org/wiki/Goran_Visnjic
Gordie Howe	http://en.wikipedia.org/wiki/Gordie_Howe
Gordon Banks	http://en.wikipedia.org/wiki/Gordon_Banks
Gordon Banks	http://en.wikipedia.org/wiki/Gordon_Banks_(politician)
Gordon Birtwistle	http://en.wikipedia.org/wiki/Gordon_Birtwistle
Gordon Brown	http://en.wikipedia.org/wiki/Gordon_Brown
Gordon Cooper	http://en.wikipedia.org/wiki/Gordon_Cooper
Gordon Douglas	http://en.wikipedia.org/wiki/Gordon_Douglas_(director)
Gordon E. Sawyer	http://en.wikipedia.org/wiki/Gordon_E._Sawyer
Gordon Getty	http://en.wikipedia.org/wiki/Gordon_Getty
Gordon Gould	http://en.wikipedia.org/wiki/Gordon_Gould
Gordon Gray	http://en.wikipedia.org/wiki/Gordon_Gray_(politician)
Gordon Henderson	http://en.wikipedia.org/wiki/Gordon_Henderson_(politician)
Gordon Hinckley	http://en.wikipedia.org/wiki/Gordon_Hinckley
Gordon Humphrey	http://en.wikipedia.org/wiki/Gordon_Humphrey
Gordon J. Humphrey	http://en.wikipedia.org/wiki/Gordon_J._Humphrey
Gordon Jackson	http://en.wikipedia.org/wiki/Gordon_Jackson_(actor)
Gordon Johncock	http://en.wikipedia.org/wiki/Gordon_Johncock
Gordon Jump	http://en.wikipedia.org/wiki/Gordon_Jump
Gordon Lightfoot	http://en.wikipedia.org/wiki/Gordon_Lightfoot
Gordon MacRae	http://en.wikipedia.org/wiki/Gordon_MacRae
Gordon Marsden	http://en.wikipedia.org/wiki/Gordon_Marsden
Gordon Moore	http://en.wikipedia.org/wiki/Gordon_Moore
Gordon Parks	http://en.wikipedia.org/wiki/Gordon_Parks
Gordon R. Dickson	http://en.wikipedia.org/wiki/Gordon_R._Dickson
Gordon R. England	http://en.wikipedia.org/wiki/Gordon_R._England
Gordon Ramsay	http://en.wikipedia.org/wiki/Gordon_Ramsay
Gordon Smith	http://en.wikipedia.org/wiki/Gordon_H._Smith
Gordon W. Allport	http://en.wikipedia.org/wiki/Gordon_W._Allport
Gordon Waller	http://en.wikipedia.org/wiki/Gordon_Waller
Gore Vidal	http://en.wikipedia.org/wiki/Gore_Vidal
Gottfried August B�rger+A5675	http://en.wikipedia.org/wiki/Gottfried_August_B%C3%BCrger
Gottfried Benn	http://en.wikipedia.org/wiki/Gottfried_Benn
Gottfried Leibniz	http://en.wikipedia.org/wiki/Gottfried_Leibniz
Gotthold Ephraim Lessing	http://en.wikipedia.org/wiki/Gotthold_Ephraim_Lessing
Gough Whitlam	http://en.wikipedia.org/wiki/Gough_Whitlam
Gouverneur Kemble Warren	http://en.wikipedia.org/wiki/Gouverneur_Kemble_Warren
Gouverneur Morris	http://en.wikipedia.org/wiki/Gouverneur_Morris
Grace Abbott	http://en.wikipedia.org/wiki/Grace_Abbott
Grace Darling	http://en.wikipedia.org/wiki/Grace_Darling
Grace Jones	http://en.wikipedia.org/wiki/Grace_Jones
Grace Kelly	http://en.wikipedia.org/wiki/Grace_Kelly
Grace Lumpkin	http://en.wikipedia.org/wiki/Grace_Lumpkin
Grace Metalious	http://en.wikipedia.org/wiki/Grace_Metalious
Grace Murray Hopper	http://en.wikipedia.org/wiki/Grace_Murray_Hopper
Grace Napolitano	http://en.wikipedia.org/wiki/Grace_Napolitano
Grace Paley	http://en.wikipedia.org/wiki/Grace_Paley
Grace Slick	http://en.wikipedia.org/wiki/Grace_Slick
Grace Zabriskie	http://en.wikipedia.org/wiki/Grace_Zabriskie
Gracie Allen	http://en.wikipedia.org/wiki/Gracie_Allen
Graeme Allwright	http://en.wikipedia.org/wiki/Graeme_Allwright
Graeme Morrice	http://en.wikipedia.org/wiki/Graeme_Morrice
Graeme Smith	http://en.wikipedia.org/wiki/Graeme_Smith
Graham Allen	http://en.wikipedia.org/wiki/Graham_Allen_(politician)
Graham Bond	http://en.wikipedia.org/wiki/Graham_Bond
Graham Brady	http://en.wikipedia.org/wiki/Graham_Brady
Graham Chapman	http://en.wikipedia.org/wiki/Graham_Chapman
Graham Coxon	http://en.wikipedia.org/wiki/Graham_Coxon
Graham Evans	http://en.wikipedia.org/wiki/Graham_Evans
Graham Greene	http://en.wikipedia.org/wiki/Graham_Greene
Graham Greene	http://en.wikipedia.org/wiki/Graham_Greene
Graham Jones	http://en.wikipedia.org/wiki/Graham_Jones_(politician)
Graham Kerr	http://en.wikipedia.org/wiki/Graham_Kerr
Graham Nash	http://en.wikipedia.org/wiki/Graham_Nash
Graham Nelson	http://en.wikipedia.org/wiki/Graham_Nelson
Graham Norton	http://en.wikipedia.org/wiki/Graham_Norton
Graham Parker	http://en.wikipedia.org/wiki/Graham_Parker
Graham Russell	http://en.wikipedia.org/wiki/Graham_Russell
Graham Stringer	http://en.wikipedia.org/wiki/Graham_Stringer
Graham Stuart	http://en.wikipedia.org/wiki/Graham_Stuart_(UK_politician)
Graham Swift	http://en.wikipedia.org/wiki/Graham_Swift
Grahame Morris	http://en.wikipedia.org/wiki/Grahame_Morris
Gram Parsons	http://en.wikipedia.org/wiki/Gram_Parsons
Grand Duke Henri	http://en.wikipedia.org/wiki/Grand_Duke_Henri
Grand Verbalizer Funkin-Lesson	http://en.wikipedia.org/wiki/X-Clan
Grandma Moses	http://en.wikipedia.org/wiki/Grandma_Moses
Grandmaster Flash	http://en.wikipedia.org/wiki/Grandmaster_Flash
Grandpa Jones	http://en.wikipedia.org/wiki/Grandpa_Jones
Grant Hill	http://en.wikipedia.org/wiki/Grant_Hill
Grant Lee Phillips	http://en.wikipedia.org/wiki/Grant_Lee_Phillips
Grant Mitchell	http://en.wikipedia.org/wiki/Grant_Mitchell_(actor)
Grant Sawyer	http://en.wikipedia.org/wiki/Grant_Sawyer
Grant Shapps	http://en.wikipedia.org/wiki/Grant_Shapps
Grant Shaud	http://en.wikipedia.org/wiki/Grant_Shaud
Grant Show	http://en.wikipedia.org/wiki/Grant_Show
Grant Tinker	http://en.wikipedia.org/wiki/Grant_Tinker
Grant Withers	http://en.wikipedia.org/wiki/Grant_Withers
Grant Wood	http://en.wikipedia.org/wiki/Grant_Wood
Granville Hicks	http://en.wikipedia.org/wiki/Granville_Hicks
Granville Sharp	http://en.wikipedia.org/wiki/Granville_Sharp
Gray Davis	http://en.wikipedia.org/wiki/Gray_Davis
Graydon Carter	http://en.wikipedia.org/wiki/Graydon_Carter
Green Gartside	http://en.wikipedia.org/wiki/Green_Gartside
Greer Garson	http://en.wikipedia.org/wiki/Greer_Garson
Greg Bear	http://en.wikipedia.org/wiki/Greg_Bear
Greg Behrendt	http://en.wikipedia.org/wiki/Greg_Behrendt
Greg Clark	http://en.wikipedia.org/wiki/Greg_Clark
Greg Evigan	http://en.wikipedia.org/wiki/Greg_Evigan
Greg Ginn	http://en.wikipedia.org/wiki/Greg_Ginn
Greg Graffin	http://en.wikipedia.org/wiki/Greg_Graffin
Greg Ham	http://en.wikipedia.org/wiki/Greg_Ham
Greg Hands	http://en.wikipedia.org/wiki/Greg_Hands
Greg Kinnear	http://en.wikipedia.org/wiki/Greg_Kinnear
Greg Knight	http://en.wikipedia.org/wiki/Greg_Knight
Greg Lake	http://en.wikipedia.org/wiki/Greg_Lake
Greg Lauren	http://en.wikipedia.org/wiki/Greg_Lauren
Greg Laurie	http://en.wikipedia.org/wiki/Greg_Laurie
Greg Lisher	http://en.wikipedia.org/wiki/Greg_Lisher
Greg Louganis	http://en.wikipedia.org/wiki/Greg_Louganis
Greg Maddux	http://en.wikipedia.org/wiki/Greg_Maddux
Greg Mankiw	http://en.wikipedia.org/wiki/Greg_Mankiw
Greg Morris	http://en.wikipedia.org/wiki/Greg_Morris
Greg Mulholland	http://en.wikipedia.org/wiki/Greg_Mulholland
Greg Norman	http://en.wikipedia.org/wiki/Greg_Norman
Greg Palast	http://en.wikipedia.org/wiki/Greg_Palast
Greg Proops	http://en.wikipedia.org/wiki/Greg_Proops
Greg Walden	http://en.wikipedia.org/wiki/Greg_Walden
Gregg Allman	http://en.wikipedia.org/wiki/Gregg_Allman
Gregg Harper	http://en.wikipedia.org/wiki/Gregg_Harper
Gregg Henry	http://en.wikipedia.org/wiki/Gregg_Henry
Gregg McClymont	http://en.wikipedia.org/wiki/Gregg_McClymont
Gregg Rolie	http://en.wikipedia.org/wiki/Gregg_Rolie
Gregor Mendel	http://en.wikipedia.org/wiki/Gregor_Mendel
Gregor Strasser	http://en.wikipedia.org/wiki/Gregor_Strasser
Gregory Barker	http://en.wikipedia.org/wiki/Gregory_Barker
Gregory Bateson	http://en.wikipedia.org/wiki/Gregory_Bateson
Gregory Baylor	http://en.wikipedia.org/wiki/Gregory_Baylor
Gregory Benford	http://en.wikipedia.org/wiki/Gregory_Benford
Gregory Breit	http://en.wikipedia.org/wiki/Gregory_Breit
Gregory Campbell	http://en.wikipedia.org/wiki/Gregory_Campbell_(politician)
Gregory Corso	http://en.wikipedia.org/wiki/Gregory_Corso
Gregory Harrison	http://en.wikipedia.org/wiki/Gregory_Harrison
Gregory Hines	http://en.wikipedia.org/wiki/Gregory_Hines
Gregory Meeks	http://en.wikipedia.org/wiki/Gregory_Meeks
Gregory Peck	http://en.wikipedia.org/wiki/Gregory_Peck
Gregory Scarpa, Sr.	http://en.wikipedia.org/wiki/Gregory_Scarpa%2C_Sr.
Gregory Smith	http://en.wikipedia.org/wiki/Gregory_Smith_(actor)
Gregory Vlastos	http://en.wikipedia.org/wiki/Gregory_Smith_(actor)
Gregory XVI	http://en.wikipedia.org/wiki/Gregory_Smith_(actor)
Gresham Barrett	http://en.wikipedia.org/wiki/Gregory_XVI
Greta Garbo	http://en.wikipedia.org/wiki/Greta_Garbo
Greta Scacchi	http://en.wikipedia.org/wiki/Greta_Scacchi
Greta Van Susteren	http://en.wikipedia.org/wiki/Greta_Van_Susteren
Gretchen Mol	http://en.wikipedia.org/wiki/Gretchen_Mol
Gretchen Wilson	http://en.wikipedia.org/wiki/Gretchen_Wilson
Griff Rhys Jones	http://en.wikipedia.org/wiki/Griff_Rhys_Jones
Griffin Dunne	http://en.wikipedia.org/wiki/Griffin_Dunne
Grinling Gibbons	http://en.wikipedia.org/wiki/Grinling_Gibbons
Groucho Marx	http://en.wikipedia.org/wiki/Groucho_Marx
Grover Cleveland	http://en.wikipedia.org/wiki/Grover_Cleveland
Grover Cleveland Alexander	http://en.wikipedia.org/wiki/Grover_Cleveland_Alexander
Grover Norquist	http://en.wikipedia.org/wiki/Grover_Norquist
Guglielmo Marconi	http://en.wikipedia.org/wiki/Guglielmo_Marconi
Guido Cavalcanti	http://en.wikipedia.org/wiki/Guido_Cavalcanti
Guido Reni	http://en.wikipedia.org/wiki/Guido_Reni
Guido van Rossum	http://en.wikipedia.org/wiki/Guido_van_Rossum
Guillaume Amontons	http://en.wikipedia.org/wiki/Guillaume_Amontons
Guillaume Apollinaire	http://en.wikipedia.org/wiki/Guillaume_Apollinaire
Guillaume Dufay	http://en.wikipedia.org/wiki/Guillaume_Dufay
Guillaume Farel	http://en.wikipedia.org/wiki/Guillaume_Farel
Guillaume Soro	http://en.wikipedia.org/wiki/Guillaume_Soro
Guillermo Cabrera Infante	http://en.wikipedia.org/wiki/Guillermo_Cabrera_Infante
Guillermo Coria	http://en.wikipedia.org/wiki/Guillermo_Coria
Guillermo del Toro	http://en.wikipedia.org/wiki/Guillermo_del_Toro
Guillermo Endara	http://en.wikipedia.org/wiki/Guillermo_Endara
Guinevere Turner	http://en.wikipedia.org/wiki/Guinevere_Turner
Gulbuddin Hekmatyar	http://en.wikipedia.org/wiki/Gulbuddin_Hekmatyar
Gulshan Grover	http://en.wikipedia.org/wiki/Gulshan_Grover
Gummo Marx	http://en.wikipedia.org/wiki/Gummo_Marx
Gunnar Gunnarsson	http://en.wikipedia.org/wiki/Gunnar_Gunnarsson
Gunnar Myrdal	http://en.wikipedia.org/wiki/Gunnar_Myrdal
G�nter Grass	http://en.wikipedia.org/wiki/G%C3%BCnter_Grass
Gunther von Hagens	http://en.wikipedia.org/wiki/Gunther_von_Hagens
G�nther von Kluge	http://en.wikipedia.org/wiki/G%C3%BCnther_von_Kluge
Gurbanguly Berdimuhamedow	http://en.wikipedia.org/wiki/Gurbanguly_Berdimuhamedow
Gus Bilirkis	http://en.wikipedia.org/wiki/Gus_Bilirkis
Gus Grissom	http://en.wikipedia.org/wiki/Gus_Grissom
Gus Savage	http://en.wikipedia.org/wiki/Gus_Savage
Gus Van Sant	http://en.wikipedia.org/wiki/Gus_Van_Sant
Gus Yatron	http://en.wikipedia.org/wiki/Gus_Yatron
Gustaf Dal�n+A5721	http://en.wikipedia.org/wiki/Gustaf_Dal%C3%A9n
Gustav Adolph the Great	http://en.wikipedia.org/wiki/Gustavus_Adolphus_of_Sweden
Gustav Bauer	http://en.wikipedia.org/wiki/Gustav_Bauer
Gustav Heinemann	http://en.wikipedia.org/wiki/Gustav_Heinemann
Gustav Hertz	http://en.wikipedia.org/wiki/Gustav_Hertz
Gustav Holst	http://en.wikipedia.org/wiki/Gustav_Holst
Gustav Klimt	http://en.wikipedia.org/wiki/Gustav_Klimt
Gustav Knuth	http://en.wikipedia.org/wiki/Gustav_Knuth
Gustav Krupp	http://en.wikipedia.org/wiki/Gustav_Krupp
Gustav Mahler	http://en.wikipedia.org/wiki/Gustav_Mahler
Gustav Robert Kirchhoff	http://en.wikipedia.org/wiki/Gustav_Robert_Kirchhoff
Gustav Stresemann	http://en.wikipedia.org/wiki/Gustav_Stresemann
Gustav V	http://en.wikipedia.org/wiki/Gustav_V
Gustave Charpentier	http://en.wikipedia.org/wiki/Gustave_Charpentier
Gustave Courbet	http://en.wikipedia.org/wiki/Gustave_Courbet
Gustave Dor�	http://en.wikipedia.org/wiki/Gustave_Dor%C3%A9
Gustave Eiffel	http://en.wikipedia.org/wiki/Gustave_Eiffel
Gustave Flaubert	http://en.wikipedia.org/wiki/Gustave_Flaubert
Guto Bebb	http://en.wikipedia.org/wiki/Guto_Bebb
Guy Berryman	http://en.wikipedia.org/wiki/Guy_Berryman
Guy Davenport	http://en.wikipedia.org/wiki/Guy_Davenport
Guy de Maupassant	http://en.wikipedia.org/wiki/Guy_de_Maupassant
Guy Fawkes	http://en.wikipedia.org/wiki/Guy_Fawkes
Guy Gavriel Kay	http://en.wikipedia.org/wiki/Guy_Gavriel_Kay
Guy Hamilton	http://en.wikipedia.org/wiki/Guy_Hamilton
Guy Kawasaki	http://en.wikipedia.org/wiki/Guy_Kawasaki
Guy Kibbee	http://en.wikipedia.org/wiki/Guy_Kibbee
Guy Liddell	http://en.wikipedia.org/wiki/Guy_Liddell
Guy Lombardo	http://en.wikipedia.org/wiki/Guy_Lombardo
Guy Madison	http://en.wikipedia.org/wiki/Guy_Madison
Guy Opperman	http://en.wikipedia.org/wiki/Guy_Opperman
Guy Pearce	http://en.wikipedia.org/wiki/Guy_Pearce
Guy Ritchie	http://en.wikipedia.org/wiki/Guy_Ritchie
Guy V. Molinari	http://en.wikipedia.org/wiki/Guy_V._Molinari
Guy Vander Jagt	http://en.wikipedia.org/wiki/Guy_Vander_Jagt
Guy Verhofstadt	http://en.wikipedia.org/wiki/Guy_Verhofstadt
Guy Verhofstadt	http://en.wikipedia.org/wiki/Guy_Verhofstadt
Guy Williams	http://en.wikipedia.org/wiki/Guy_Williams
Gwen Ifill	http://en.wikipedia.org/wiki/Gwen_Ifill
Gwen Moore	http://en.wikipedia.org/wiki/Gwen_Moore
Gwen Stefani	http://en.wikipedia.org/wiki/Gwen_Stefani
Gwen Verdon	http://en.wikipedia.org/wiki/Gwen_Verdon
Gwendolyn Bennett	http://en.wikipedia.org/wiki/Gwendolyn_Bennett
Gwendolyn Brooks	http://en.wikipedia.org/wiki/Gwendolyn_Brooks
Gwendolyn MacEwen	http://en.wikipedia.org/wiki/Gwendolyn_MacEwen
Gwyneth Paltrow	http://en.wikipedia.org/wiki/Gwyneth_Paltrow
Gyanendra Bir Bikram Shah Dev	http://en.wikipedia.org/wiki/Gyanendra_Bir_Bikram_Shah_Dev
Gy�rgy Ligeti Ligeti	http://en.wikipedia.org/wiki/Gy%C3%B6rgy_Ligeti
Gypsy Abbott	http://en.wikipedia.org/wiki/Gypsy_Abbott
Gypsy Rose Lee	http://en.wikipedia.org/wiki/Gypsy_Rose_Lee
Gyude Bryant	http://en.wikipedia.org/wiki/Gyude_Bryant
Gyula Horn	http://en.wikipedia.org/wiki/Gyula_Horn
H. Bruce Humberstone	http://en.wikipedia.org/wiki/H._Bruce_Humberstone
H. D.	http://en.wikipedia.org/wiki/H._D.
H. E. Bates	http://en.wikipedia.org/wiki/H._E._Bates
H. G. Wells	http://en.wikipedia.org/wiki/H._G._Wells
H. H. Holmes	http://en.wikipedia.org/wiki/H._H._Holmes
H. H. Munro	http://en.wikipedia.org/wiki/H._H._Munro
H. James Saxton	http://en.wikipedia.org/wiki/H._James_Saxton
H. L. Davis	http://en.wikipedia.org/wiki/H._L._Davis
H. L. Hunt	http://en.wikipedia.org/wiki/H._L._Hunt
H. L. Mencken	http://en.wikipedia.org/wiki/H._L._Mencken
H. Lee Scott	http://en.wikipedia.org/wiki/H._Lee_Scott
H. Lee Scott Jr.	http://en.wikipedia.org/wiki/H._Lee_Scott_Jr.
H. P. Blavatsky	http://en.wikipedia.org/wiki/H._P._Blavatsky
H. P. Lovecraft	http://en.wikipedia.org/wiki/H._P._Lovecraft
H. R. Giger	http://en.wikipedia.org/wiki/H._R._Giger
H. R. Haldeman	http://en.wikipedia.org/wiki/H._R._Haldeman
H. Rap Brown	http://en.wikipedia.org/wiki/H._Rap_Brown
H. Rider Haggard	http://en.wikipedia.org/wiki/H._Rider_Haggard
H. Ross Perot	http://en.wikipedia.org/wiki/H._Ross_Perot
H. Wayne Huizenga	http://en.wikipedia.org/wiki/H._Wayne_Huizenga
Haakon I Adalsteinsfostre	http://en.wikipedia.org/wiki/Haakon_I_Adalsteinsfostre
Haakon IV Haakonsson	http://en.wikipedia.org/wiki/Haakon_IV_Haakonsson
Hack Wilson	http://en.wikipedia.org/wiki/Hack_Wilson
Hadassah Lieberman	http://en.wikipedia.org/wiki/Hadassah_Lieberman
Hafez al-Assad	http://en.wikipedia.org/wiki/Hafez_al-Assad
Hafizullah Amin	http://en.wikipedia.org/wiki/Hafizullah_Amin
Haifa Wehbe	http://en.wikipedia.org/wiki/Haifa_Wehbe
Haile Selassie	http://en.wikipedia.org/wiki/Haile_Selassie
Haing S. Ngor	http://en.wikipedia.org/wiki/Haing_S._Ngor
Hakeem Abdul-Samad	http://en.wikipedia.org/wiki/The_Boys_%28band%29
Hakeem Olajuwon	http://en.wikipedia.org/wiki/Hakeem_Olajuwon
Haki R. Madhubuti	http://en.wikipedia.org/wiki/Haki_R._Madhubuti
Hal Ashby	http://en.wikipedia.org/wiki/Hal_Ashby
Hal Daub	http://en.wikipedia.org/wiki/Hal_Daub
Hal Hartley	http://en.wikipedia.org/wiki/Hal_Hartley
Hal Holbrook	http://en.wikipedia.org/wiki/Hal_Holbrook
Hal Linden	http://en.wikipedia.org/wiki/Hal_Linden
Hal Lindsey	http://en.wikipedia.org/wiki/Hal_Lindsey
Hal Roach	http://en.wikipedia.org/wiki/Hal_Roach
Hal Rogers	http://en.wikipedia.org/wiki/Hal_Rogers
Hal Sparks	http://en.wikipedia.org/wiki/Hal_Sparks
Hale Boggs	http://en.wikipedia.org/wiki/Hale_Boggs
Haley Barbour	http://en.wikipedia.org/wiki/Haley_Barbour
Haley Barbour	http://en.wikipedia.org/wiki/Haley_Barbour
Haley Joel Osment	http://en.wikipedia.org/wiki/Haley_Joel_Osment
Halld�r �sgr�msson	http://en.wikipedia.org/wiki/Halld%C3%B3r_%C3%81sgr%C3%Admsson
Halle Berry	http://en.wikipedia.org/wiki/Halle_Berry
Ham Lini	http://en.wikipedia.org/wiki/Ham_Lini
Hama Amadou	http://en.wikipedia.org/wiki/Hama_Amadou
Hamad bin Isa Al Khalifa	http://en.wikipedia.org/wiki/Hamad_bin_Isa_Al_Khalifa
Hamad bin Jassim bin Jaber Al Thani	http://en.wikipedia.org/wiki/Hamad_bin_Jassim_bin_Jaber_Al_Thani
Hamad bin Khalifa Al Thani	http://en.wikipedia.org/wiki/Hamad_bin_Khalifa_Al_Thani
Hamid Karzai	http://en.wikipedia.org/wiki/Hamid_Karzai
Hamid Karzai	http://en.wikipedia.org/wiki/Hamid_Karzai
Hamilton Fish	http://en.wikipedia.org/wiki/Hamilton_Fish
Hamilton Fish, Jr.	http://en.wikipedia.org/wiki/Hamilton_Fish
Hamilton Jordan	http://en.wikipedia.org/wiki/Hamilton_Jordan
Hamlin Garland	http://en.wikipedia.org/wiki/Hamlin_Garland
Han Duck Soo	http://en.wikipedia.org/wiki/Han_Duck_Soo
Han Myung Sook	http://en.wikipedia.org/wiki/Han_Myung_Sook
Hank Aaron	http://en.wikipedia.org/wiki/Hank_Aaron
Hank Azaria	http://en.wikipedia.org/wiki/Hank_Azaria
Hank Ballard	http://en.wikipedia.org/wiki/Hank_Ballard
Hank Brown	http://en.wikipedia.org/wiki/Hank_Brown
Hank Brown	http://en.wikipedia.org/wiki/Hank_Brown
Hank Garland	http://en.wikipedia.org/wiki/Hank_Garland
Hank Greenberg	http://en.wikipedia.org/wiki/Hank_Greenberg
Hank Johnson	http://en.wikipedia.org/wiki/Hank_Johnson
Hank Jones	http://en.wikipedia.org/wiki/Hank_Jones
Hank Ketcham	http://en.wikipedia.org/wiki/Hank_Ketcham
Hank Mann	http://en.wikipedia.org/wiki/Hank_Mann
Hank Penny	http://en.wikipedia.org/wiki/Hank_Penny
Hank Stram	http://en.wikipedia.org/wiki/Hank_Stram
Hank Williams III	http://en.wikipedia.org/wiki/Hank_Williams_III
Hank Williams, Jr.	http://en.wikipedia.org/wiki/Hank_Williams%2C_Jr.
Hank Williams, Sr.	http://en.wikipedia.org/wiki/Hank_Williams%2C_Sr.
Hannah Arendt	http://en.wikipedia.org/wiki/Hannah_Arendt
Hannes Alfv�n	http://en.wikipedia.org/wiki/Hannes_Alfv%C3%A9n
Hannibal Hamlin	http://en.wikipedia.org/wiki/Hannibal_Hamlin
Hanoi Hannah	http://en.wikipedia.org/wiki/Hanoi_Hannah
Hans Adam II	http://en.wikipedia.org/wiki/Hans_Adam_II
Hans Alfredson	http://en.wikipedia.org/wiki/Hans_Alfredson
Hans Bethe	http://en.wikipedia.org/wiki/Hans_Bethe
Hans Blix	http://en.wikipedia.org/wiki/Hans_Blix
Hans Burgkmair	http://en.wikipedia.org/wiki/Hans_Burgkmair
Hans Christian Andersen	http://en.wikipedia.org/wiki/Hans_Christian_Andersen
Hans Christian Oersted	http://en.wikipedia.org/wiki/Hans_Christian_Oersted
Hans Daniel Hassenpflug	http://en.wikipedia.org/wiki/Hans_Daniel_Hassenpflug
Hans Enoksen	http://en.wikipedia.org/wiki/Hans_Enoksen
Hans Filbinger	http://en.wikipedia.org/wiki/Hans_Filbinger
Hans Fischer	http://en.wikipedia.org/wiki/Hans_Fischer
Hans Frank	http://en.wikipedia.org/wiki/Hans_Frank
Hans Fritzsche	http://en.wikipedia.org/wiki/Hans_Fritzsche
Hans G. Dehmelt	http://en.wikipedia.org/wiki/Hans_G._Dehmelt
Hans Geiger	http://en.wikipedia.org/wiki/Hans_Geiger
Hans Heinrich Lammers	http://en.wikipedia.org/wiki/Hans_Heinrich_Lammers
Hans Holbein the Elder	http://en.wikipedia.org/wiki/Hans_Holbein_the_Elder
Hans Holbein the Younger	http://en.wikipedia.org/wiki/Hans_Holbein_the_Younger
Hans Luther	http://en.wikipedia.org/wiki/Hans_Luther
Hans Memling	http://en.wikipedia.org/wiki/Hans_Memling
Hans Speidel	http://en.wikipedia.org/wiki/Hans_Speidel
Hans Svane	http://en.wikipedia.org/wiki/Hans_Svane
Hans Tausen	http://en.wikipedia.org/wiki/Hans_Tausen
Hans von Euler-Chelpin	http://en.wikipedia.org/wiki/Hans_von_Euler-Chelpin
Hans Werner Henze	http://en.wikipedia.org/wiki/Hans_Werner_Henze
Hans Zimmer	http://en.wikipedia.org/wiki/Hans_Zimmer
Hans-Georg Gadamer	http://en.wikipedia.org/wiki/Hans-Georg_Gadamer
Hany Abu-Assad	http://en.wikipedia.org/wiki/Hany_Abu-Assad
Har Mar Superstar	http://en.wikipedia.org/wiki/Har_Mar_Superstar
Harald I	http://en.wikipedia.org/wiki/Harald_I
Harald III	http://en.wikipedia.org/wiki/Harald_III_of_Norway
Harald IV	http://en.wikipedia.org/wiki/Harald_IV
Harald V	http://en.wikipedia.org/wiki/Harald_V
Hardy Amies	http://en.wikipedia.org/wiki/Hardy_Amies
Harlan Cleveland	http://en.wikipedia.org/wiki/Harlan_Cleveland
Harlan Ellison	http://en.wikipedia.org/wiki/Harlan_Ellison
Harlan Fiske Stone	http://en.wikipedia.org/wiki/Harlan_Fiske_Stone
Harley O. Staggers, Jr.	http://en.wikipedia.org/wiki/Harley_O._Staggers%2C_Jr.
Harmon Killebrew	http://en.wikipedia.org/wiki/Harmon_Killebrew
Harmony Korine	http://en.wikipedia.org/wiki/Harmony_Korine
Harold Alfond	http://en.wikipedia.org/wiki/Harold_Alfond
Harold Arlen	http://en.wikipedia.org/wiki/Harold_Arlen
Harold Becker	http://en.wikipedia.org/wiki/Harold_Becker
Harold Bell Wright	http://en.wikipedia.org/wiki/Harold_Bell_Wright
Harold Bloom	http://en.wikipedia.org/wiki/Harold_Bloom
Harold Brodkey	http://en.wikipedia.org/wiki/Harold_Brodkey
Harold Brown	http://en.wikipedia.org/wiki/Harold_Brown_(Secretary_of_Defense)
Harold Budd	http://en.wikipedia.org/wiki/Harold_Budd
Harold C. Urey	http://en.wikipedia.org/wiki/Harold_C._Urey
Harold E. Ford, Jr.	http://en.wikipedia.org/wiki/Harold_E._Ford%2C_Jr.
Harold Ford	http://en.wikipedia.org/wiki/Harold_Ford
Harold Ford, Sr.	http://en.wikipedia.org/wiki/Harold_Ford%2C_Sr.
Harold Gould	http://en.wikipedia.org/wiki/Harold_Gould
Harold Harefoot	http://en.wikipedia.org/wiki/Harold_Harefoot
Harold Hunter	http://en.wikipedia.org/wiki/Harold_Hunter
Harold Ickes	http://en.wikipedia.org/wiki/Harold_L._Ickes
Harold L. Volkmer	http://en.wikipedia.org/wiki/Harold_L._Volkmer
Harold Lloyd	http://en.wikipedia.org/wiki/Harold_Lloyd
Harold Macmillan	http://en.wikipedia.org/wiki/Harold_Macmillan
Harold McGee	http://en.wikipedia.org/wiki/Harold_McGee
Harold Nicholas	http://en.wikipedia.org/wiki/Harold_Nicholas
Harold Perrineau, Jr.	http://en.wikipedia.org/wiki/Harold_Perrineau%2C_Jr.
Harold Pinter	http://en.wikipedia.org/wiki/Harold_Pinter
Harold Ramis	http://en.wikipedia.org/wiki/Harold_Ramis
Harold Robbins	http://en.wikipedia.org/wiki/Harold_Robbins
Harold Rogers	http://en.wikipedia.org/wiki/Hal_Rogers
Harold Russell	http://en.wikipedia.org/wiki/Harold_Russell
Harold Shipman	http://en.wikipedia.org/wiki/Harold_Shipman
Harold Stassen	http://en.wikipedia.org/wiki/Harold_Stassen
Harold W. McGraw III	http://en.wikipedia.org/wiki/Harold_W._McGraw_III
Harold W. Ross	http://en.wikipedia.org/wiki/Harold_W._Ross
Harold Washington	http://en.wikipedia.org/wiki/Harold_Washington
Harold Wilson	http://en.wikipedia.org/wiki/Harold_Wilson
Harper Lee	http://en.wikipedia.org/wiki/Harper_Lee
Harpo Marx	http://en.wikipedia.org/wiki/Harpo_Marx
Harriet Ann Jacobs	http://en.wikipedia.org/wiki/Harriet_Ann_Jacobs
Harriet Beecher Stowe	http://en.wikipedia.org/wiki/Harriet_Beecher_Stowe
Harriet E. Wilson	http://en.wikipedia.org/wiki/Harriet_E._Wilson
Harriet Goodhue Hosmer	http://en.wikipedia.org/wiki/Harriet_Goodhue_Hosmer
Harriet Harman	http://en.wikipedia.org/wiki/Harriet_Harman
Harriet Hilliard	http://en.wikipedia.org/wiki/Harriet_Hilliard
Harriet MacGibbon	http://en.wikipedia.org/wiki/Harriet_MacGibbon
Harriet Martineau	http://en.wikipedia.org/wiki/Harriet_Martineau
Harriet Miers	http://en.wikipedia.org/wiki/Harriet_Miers
Harriet Monroe	http://en.wikipedia.org/wiki/Harriet_Monroe
Harriet Tubman	http://en.wikipedia.org/wiki/Harriet_Tubman
Harriett Baldwin	http://en.wikipedia.org/wiki/Harriett_Baldwin
Harris W. Fawell	http://en.wikipedia.org/wiki/Harris_W._Fawell
Harris Wofford	http://en.wikipedia.org/wiki/Harris_Wofford
Harrison Ford	http://en.wikipedia.org/wiki/Harrison_Ford
Harrison Page	http://en.wikipedia.org/wiki/Harrison_Page
Harry Anderson	http://en.wikipedia.org/wiki/Harry_Anderson
Harry Andrews	http://en.wikipedia.org/wiki/Harry_Andrews
Harry Babbitt	http://en.wikipedia.org/wiki/Harry_Babbitt
Harry Beck	http://en.wikipedia.org/wiki/Harry_Beck
Harry Belafonte	http://en.wikipedia.org/wiki/Harry_Belafonte
Harry Blackmun	http://en.wikipedia.org/wiki/Harry_Blackmun
Harry Browne	http://en.wikipedia.org/wiki/Harry_Browne
Harry Carey, Jr.	http://en.wikipedia.org/wiki/Harry_Carey%2C_Jr.
Harry Carey, Sr.	http://en.wikipedia.org/wiki/Harry_Carey_%28actor_born_1878%29
Harry Chapin	http://en.wikipedia.org/wiki/Harry_Chapin
Harry Connick, Jr.	http://en.wikipedia.org/wiki/Harry_Connick%2C_Jr.
Harry Dean Stanton	http://en.wikipedia.org/wiki/Harry_Dean_Stanton
Harry F. Byrd	http://en.wikipedia.org/wiki/Harry_F._Byrd
Harry F. Byrd, Jr.	http://en.wikipedia.org/wiki/Harry_F._Byrd%2C_Jr.
Harry Goz	http://en.wikipedia.org/wiki/Harry_Goz
Harry Hamlin	http://en.wikipedia.org/wiki/Harry_Hamlin
Harry Harrison	http://en.wikipedia.org/wiki/Harry_Harrison
Harry Hay	http://en.wikipedia.org/wiki/Harry_Hay
Harry Houdini	http://en.wikipedia.org/wiki/Harry_Houdini
Harry James	http://en.wikipedia.org/wiki/Harry_James
Harry Knowles	http://en.wikipedia.org/wiki/Harry_Knowles
Harry Langdon	http://en.wikipedia.org/wiki/Harry_Langdon
Harry Leon Wilson	http://en.wikipedia.org/wiki/Harry_Leon_Wilson
Harry Lloyd Hopkins	http://en.wikipedia.org/wiki/Harry_Lloyd_Hopkins
Harry Mark Petrakis	http://en.wikipedia.org/wiki/Harry_Mark_Petrakis
Harry Mitchell	http://en.wikipedia.org/wiki/Harry_Mitchell
Harry Morgan	http://en.wikipedia.org/wiki/Harry_Morgan
Harry Nilsson	http://en.wikipedia.org/wiki/Harry_Nilsson
Harry Partch	http://en.wikipedia.org/wiki/Harry_Partch
Harry Reasoner	http://en.wikipedia.org/wiki/Harry_Reasoner
Harry Redknapp	http://en.wikipedia.org/wiki/Harry_Redknapp
Harry Reid	http://en.wikipedia.org/wiki/Harry_Reid
Harry S. Truman	http://en.wikipedia.org/wiki/Harry_S._Truman
Harry Shannon	http://en.wikipedia.org/wiki/Harry_Shannon
Harry Shearer	http://en.wikipedia.org/wiki/Harry_Shearer
Harry Simeone	http://en.wikipedia.org/wiki/Harry_Simeone
Harry Smith	http://en.wikipedia.org/wiki/Harry_Everett_Smith
Harry Stonecipher	http://en.wikipedia.org/wiki/Harry_Stonecipher
Harry Teague	http://en.wikipedia.org/wiki/Harry_Teague
Harry Vardon	http://en.wikipedia.org/wiki/Harry_Vardon
Harry von Zell	http://en.wikipedia.org/wiki/Harry_von_Zell
Harry Whittington	http://en.wikipedia.org/wiki/Harry_Whittington
Hart Bochner	http://en.wikipedia.org/wiki/Hart_Bochner
Hart Crane	http://en.wikipedia.org/wiki/Hart_Crane
Hartmann von Aue	http://en.wikipedia.org/wiki/Hartmann_von_Aue
Hartmut Michel	http://en.wikipedia.org/wiki/Hartmut_Michel
Haruki Murakami	http://en.wikipedia.org/wiki/Haruki_Murakami
Harumi Kurihara	http://en.wikipedia.org/wiki/Harumi_Kurihara
Harun al-Rashid	http://en.wikipedia.org/wiki/Harun_al-Rashid
Harvey Carignan	http://en.wikipedia.org/wiki/Harvey_Carignan
Harvey Fierstein	http://en.wikipedia.org/wiki/Harvey_Fierstein
Harvey Firestone	http://en.wikipedia.org/wiki/Harvey_Firestone
Harvey Keitel	http://en.wikipedia.org/wiki/Harvey_Keitel
Harvey Korman	http://en.wikipedia.org/wiki/Harvey_Korman
Harvey Kurtzman	http://en.wikipedia.org/wiki/Harvey_Kurtzman
Harvey Milk	http://en.wikipedia.org/wiki/Harvey_Milk
Harvey Pekar	http://en.wikipedia.org/wiki/Harvey_Pekar
Harvey Pitt	http://en.wikipedia.org/wiki/Harvey_Pitt
Harvey Weinstein	http://en.wikipedia.org/wiki/Harvey_Weinstein
Hashim Thaçi	http://en.wikipedia.org/wiki/Hashim_Tha%C3%A7i
Hasil Adkins	http://en.wikipedia.org/wiki/Hasil_Adkins
Hassan Nasrallah	http://en.wikipedia.org/wiki/Hassan_Nasrallah
Hassanal Bolkiah	http://en.wikipedia.org/wiki/Hassanal_Bolkiah
Hattie Jacques	http://en.wikipedia.org/wiki/Hattie_Jacques
Hattie McDaniel	http://en.wikipedia.org/wiki/Hattie_McDaniel
Hauk Aabel	http://en.wikipedia.org/wiki/Hauk_Aabel
Hava Alberstein	http://en.wikipedia.org/wiki/Hava_Alberstein
Havelock Ellis	http://en.wikipedia.org/wiki/Havelock_Ellis
Hayao Miyazaki	http://en.wikipedia.org/wiki/Hayao_Miyazaki
Hayden Carruth	http://en.wikipedia.org/wiki/Hayden_Carruth
Hayden Christensen	http://en.wikipedia.org/wiki/Hayden_Christensen
Hayden Fry	http://en.wikipedia.org/wiki/Hayden_Fry
Hayden Panettiere	http://en.wikipedia.org/wiki/Hayden_Panettiere
Hayley Mills	http://en.wikipedia.org/wiki/Hayley_Mills
Haylie Duff	http://en.wikipedia.org/wiki/Haylie_Duff
Hayyim Nahman Bialik	http://en.wikipedia.org/wiki/Hayyim_Nahman_Bialik
Hazel Blears	http://en.wikipedia.org/wiki/Hazel_Blears
Hazel O'Leary	http://en.wikipedia.org/wiki/Hazel_O%27Leary
Heath Ledger	http://en.wikipedia.org/wiki/Heath_Ledger
Heath Shuler	http://en.wikipedia.org/wiki/Heath_Shuler
Heather Donahue	http://en.wikipedia.org/wiki/Heather_Donahue
Heather Graham	http://en.wikipedia.org/wiki/Heather_Graham_(actress)
Heather Lauren Olson	http://en.wikipedia.org/wiki/Heather_Lauren_Olson
Heather Locklear	http://en.wikipedia.org/wiki/Heather_Locklear
Heather Mac Donald	http://en.wikipedia.org/wiki/Heather_Mac_Donald
Heather Matarazzo	http://en.wikipedia.org/wiki/Heather_Matarazzo
Heather Mills	http://en.wikipedia.org/wiki/Heather_Mills
Heather O'Rourke	http://en.wikipedia.org/wiki/Heather_O%27Rourke
Heather Small	http://en.wikipedia.org/wiki/Heather_Small
Heather Thomas	http://en.wikipedia.org/wiki/Heather_Thomas
Heather Wheeler	http://en.wikipedia.org/wiki/Heather_Wheeler
Heather Wilson	http://en.wikipedia.org/wiki/Heather_Wilson
Hecataeus of Miletus	http://en.wikipedia.org/wiki/Hecataeus_of_Miletus
Hector Berlioz	http://en.wikipedia.org/wiki/Hector_Berlioz
Hector Elizondo	http://en.wikipedia.org/wiki/Hector_Elizondo
Hector Zazou	http://en.wikipedia.org/wiki/Hector_Zazou
Hedda Hopper	http://en.wikipedia.org/wiki/Hedda_Hopper
Hedy Lamarr	http://en.wikipedia.org/wiki/Hedy_Lamarr
Hedy Lamarr	http://en.wikipedia.org/wiki/Hedy_Lamarr
Heidi Alexander	http://en.wikipedia.org/wiki/Heidi_Alexander
Heidi Fleiss	http://en.wikipedia.org/wiki/Heidi_Fleiss
Heidi Julavits	http://en.wikipedia.org/wiki/Heidi_Julavits
Heidi Klum	http://en.wikipedia.org/wiki/Heidi_Klum
Heike Kamerlingh Onnes	http://en.wikipedia.org/wiki/Heike_Kamerlingh_Onnes
Heike Makatsch	http://en.wikipedia.org/wiki/Heike_Makatsch
Heinrich Anton de Bary	http://en.wikipedia.org/wiki/Heinrich_Anton_de_Bary
Heinrich B�ll	http://en.wikipedia.org/wiki/Heinrich_B%C3%B6ll
Heinrich Bruening	http://en.wikipedia.org/wiki/Heinrich_Bruening
Heinrich Bullinger	http://en.wikipedia.org/wiki/Heinrich_Bullinger
Heinrich Harrer	http://en.wikipedia.org/wiki/Heinrich_Harrer
Heinrich Heine	http://en.wikipedia.org/wiki/Heinrich_Heine
Heinrich Hertz	http://en.wikipedia.org/wiki/Heinrich_Hertz
Heinrich Himmler	http://en.wikipedia.org/wiki/Heinrich_Himmler
Heinrich L�bke	http://en.wikipedia.org/wiki/Heinrich_L%C3%Bcbke
Heinrich Rohrer	http://en.wikipedia.org/wiki/Heinrich_Rohrer
Heinrich Schliemann	http://en.wikipedia.org/wiki/Heinrich_Schliemann
Heinrich Suso	http://en.wikipedia.org/wiki/Heinrich_Suso
Heinrich Wieland	http://en.wikipedia.org/wiki/Heinrich_Wieland
Heinz C. Prechter	http://en.wikipedia.org/wiki/Heinz_Prechter
Heinz Fischer	http://en.wikipedia.org/wiki/Heinz_Fischer
Heinz Guderian	http://en.wikipedia.org/wiki/Heinz_Guderian
Heitor Villa-Lobos	http://en.wikipedia.org/wiki/Heitor_Villa-Lobos
Helen Chenoweth-Hage	http://en.wikipedia.org/wiki/Helen_Chenoweth-Hage
Helen Clark	http://en.wikipedia.org/wiki/Helen_Clark
Helen Clark	http://en.wikipedia.org/wiki/Helen_Clark
Helen Delich Bentley	http://en.wikipedia.org/wiki/Helen_Delich_Bentley
Helen Fielding	http://en.wikipedia.org/wiki/Helen_Fielding
Helen Gallagher	http://en.wikipedia.org/wiki/Helen_Gallagher
Helen Garner	http://en.wikipedia.org/wiki/Helen_Garner
Helen Goodman	http://en.wikipedia.org/wiki/Helen_Goodman
Helen Grant	http://en.wikipedia.org/wiki/Helen_Grant_(politician)
Helen Gurley Brown	http://en.wikipedia.org/wiki/Helen_Gurley_Brown
Helen Hayes	http://en.wikipedia.org/wiki/Helen_Hayes
Helen Hokinson	http://en.wikipedia.org/wiki/Helen_Hokinson
Helen Hunt	http://en.wikipedia.org/wiki/Helen_Hunt
Helen Hunt Jackson	http://en.wikipedia.org/wiki/Helen_Hunt_Jackson
Helen Jones	http://en.wikipedia.org/wiki/Helen_Jones
Helen Keller	http://en.wikipedia.org/wiki/Helen_Keller
Helen Mirren	http://en.wikipedia.org/wiki/Helen_Mirren
Helen Reddy	http://en.wikipedia.org/wiki/Helen_Reddy
Helen Robson Walton	http://en.wikipedia.org/wiki/Helen_Robson_Walton
Helen Slater	http://en.wikipedia.org/wiki/Helen_Slater
Helen Thomas	http://en.wikipedia.org/wiki/Helen_Thomas
Helen Tucker	http://en.wikipedia.org/wiki/Helen_Tucker
Helen Vendler	http://en.wikipedia.org/wiki/Helen_Vendler
Helena Bonham Carter	http://en.wikipedia.org/wiki/Helena_Bonham_Carter
Helena Christensen	http://en.wikipedia.org/wiki/Helena_Christensen
Helene Weigel	http://en.wikipedia.org/wiki/Helene_Weigel
Hellanicus of Lesbos	http://en.wikipedia.org/wiki/Hellanicus_of_Lesbos
Helmut Berger	http://en.wikipedia.org/wiki/Helmut_Berger
Helmut Kohl	http://en.wikipedia.org/wiki/Helmut_Kohl
Helmut Lang	http://en.wikipedia.org/wiki/Helmut_Lang_(fashion_designer)
Helmut Newton	http://en.wikipedia.org/wiki/Helmut_Newton
Helmut Schmidt	http://en.wikipedia.org/wiki/Helmut_Schmidt
Helmuth von Moltke	http://en.wikipedia.org/wiki/Helmuth_James_Graf_von_Moltke
Hendrik Lorentz	http://en.wikipedia.org/wiki/Hendrik_Lorentz
Hendrik Willem van Loon	http://en.wikipedia.org/wiki/Hendrik_Willem_van_Loon
Henny Youngman	http://en.wikipedia.org/wiki/Henny_Youngman
Henri Becquerel	http://en.wikipedia.org/wiki/Henri_Becquerel
Henri Bergson	http://en.wikipedia.org/wiki/Henri_Bergson
Henri Cartier-Bresson	http://en.wikipedia.org/wiki/Henri_Cartier-Bresson
Henri de la Tour d'Auvergne	http://en.wikipedia.org/wiki/Henri_de_la_Tour_d%27Auvergne
Henri de Saint-Simon	http://en.wikipedia.org/wiki/Henri_de_Saint-Simon
Henri de Toulouse-Lautrec	http://en.wikipedia.org/wiki/Henri_de_Toulouse-Lautrec
Henri Fantin-Latour	http://en.wikipedia.org/wiki/Henri_Fantin-Latour
Henri I	http://en.wikipedia.org/wiki/Henri_I_de_Savoie,_Duc_de_Nemours
Henri II	http://en.wikipedia.org/wiki/Henry_II_of_France
Henri III	http://en.wikipedia.org/wiki/Henri_III
Henri IV	http://en.wikipedia.org/wiki/Henri_IV
Henri La Fontaine	http://en.wikipedia.org/wiki/Henri_La_Fontaine
Henri Landru	http://en.wikipedia.org/wiki/Henri_Landru
Henri Matisse	http://en.wikipedia.org/wiki/Henri_Matisse
Henri Moissan	http://en.wikipedia.org/wiki/Henri_Moissan
Henri Poincar�	http://en.wikipedia.org/wiki/Henri_Poincar%C3%A9
Henri Rousseau	http://en.wikipedia.org/wiki/Henri_Rousseau
Henri, Comte de Chambord	http://en.wikipedia.org/wiki/Henri%2C_Comte_de_Chambord
Henrietta Anne Stuart	http://en.wikipedia.org/wiki/Henrietta_Anne_Stuart
Henri-Fr�d�ric Amiel	http://en.wikipedia.org/wiki/Henri_Fr%C3%A9d%C3%A9ric_Amiel
Henrik Ibsen	http://en.wikipedia.org/wiki/Henrik_Ibsen
Henrik Tikkanen	http://en.wikipedia.org/wiki/Henrik_Tikkanen
Henri-Victor Regnault	http://en.wikipedia.org/wiki/Henri-Victor_Regnault
Henry "Scoop" Jackson	http://en.wikipedia.org/wiki/Henry_%22Scoop%22_Jackson
Henry A. Wallace	http://en.wikipedia.org/wiki/Henry_A._Wallace
Henry A. Waxman	http://en.wikipedia.org/wiki/Henry_A._Waxman
Henry Adams	http://en.wikipedia.org/wiki/Henry_Adams
Henry Addington	http://en.wikipedia.org/wiki/Henry_Addington
Henry Ainley	http://en.wikipedia.org/wiki/Henry_Ainley
Henry Armetta	http://en.wikipedia.org/wiki/Henry_Armetta
Henry Augustus Rowland	http://en.wikipedia.org/wiki/Henry_Augustus_Rowland
Henry B. Gonzalez	http://en.wikipedia.org/wiki/Henry_B._Gonzalez
Henry B. Gonzalez	http://en.wikipedia.org/wiki/Henry_B._Gonzalez
Henry B. Schacht	http://en.wikipedia.org/wiki/Henry_B._Schacht
Henry Baldwin	http://en.wikipedia.org/wiki/Henry_Baldwin_(judge)
Henry Bellingham	http://en.wikipedia.org/wiki/Henry_Bellingham_(politician)
Henry Bessemer	http://en.wikipedia.org/wiki/Henry_Bessemer
Henry Bonilla	http://en.wikipedia.org/wiki/Henry_Bonilla
Henry Box Brown	http://en.wikipedia.org/wiki/Henry_Box_Brown
Henry Brown	http://en.wikipedia.org/wiki/Henry_E._Brown,_Jr.
Henry Burghersh	http://en.wikipedia.org/wiki/Henry_Burghersh
Henry C. Carey	http://en.wikipedia.org/wiki/Henry_C._Carey
Henry Cabot Lodge	http://en.wikipedia.org/wiki/Henry_Cabot_Lodge
Henry Cabot Lodge, Jr.	http://en.wikipedia.org/wiki/Henry_Cabot_Lodge%2C_Jr.
Henry Campbell-Bannerman	http://en.wikipedia.org/wiki/Henry_Campbell-Bannerman
Henry Carter Adams	http://en.wikipedia.org/wiki/Henry_Carter_Adams
Henry Cavendish	http://en.wikipedia.org/wiki/Henry_Cavendish
Henry Cisneros	http://en.wikipedia.org/wiki/Henry_Cisneros
Henry Clay	http://en.wikipedia.org/wiki/Henry_Clay
Henry Cowell	http://en.wikipedia.org/wiki/Henry_Cowell
Henry Cuellar	http://en.wikipedia.org/wiki/Henry_Cuellar
Henry Darrow	http://en.wikipedia.org/wiki/Henry_Darrow
Henry David Thoreau	http://en.wikipedia.org/wiki/Henry_David_Thoreau
Henry de Bracton	http://en.wikipedia.org/wiki/Henry_de_Bracton
Henry de la Beche	http://en.wikipedia.org/wiki/Henry_de_la_Beche
Henry Dreyfuss	http://en.wikipedia.org/wiki/Henry_Dreyfuss
Henry Dunant	http://en.wikipedia.org/wiki/Henry_Dunant
Henry Fielding	http://en.wikipedia.org/wiki/Henry_Fielding
Henry Flynt	http://en.wikipedia.org/wiki/Henry_Flynt
Henry Fonda	http://en.wikipedia.org/wiki/Henry_Fonda
Henry Ford	http://en.wikipedia.org/wiki/Henry_Ford
Henry Ford II	http://en.wikipedia.org/wiki/Henry_Ford_II
Henry George	http://en.wikipedia.org/wiki/Henry_George
Henry Gibson	http://en.wikipedia.org/wiki/Henry_Gibson
Henry Grattan	http://en.wikipedia.org/wiki/Henry_Grattan
Henry Gwyn Jeffreys Moseley	http://en.wikipedia.org/wiki/Henry_Gwyn_Jeffreys_Moseley
Henry Hallam	http://en.wikipedia.org/wiki/Henry_Hallam
Henry Hardinge	http://en.wikipedia.org/wiki/Henry_Hardinge
Henry Harland	http://en.wikipedia.org/wiki/Henry_Harland
Henry Hathaway	http://en.wikipedia.org/wiki/Henry_Hathaway
Henry Heimlich	http://en.wikipedia.org/wiki/Henry_Heimlich
Henry Hill	http://en.wikipedia.org/wiki/Henry_Hill
Henry Hudson	http://en.wikipedia.org/wiki/Henry_Hudson
Henry Hyde	http://en.wikipedia.org/wiki/Henry_Hyde
Henry Ireton	http://en.wikipedia.org/wiki/Henry_Ireton
Henry J. Heinz	http://en.wikipedia.org/wiki/Henry_J._Heinz
Henry J. Hyde	http://en.wikipedia.org/wiki/Henry_J._Hyde
Henry J. Kaiser	http://en.wikipedia.org/wiki/Henry_J._Kaiser
Henry J. Nowak	http://en.wikipedia.org/wiki/Henry_J._Nowak
Henry James	http://en.wikipedia.org/wiki/Henry_James
Henry King	http://en.wikipedia.org/wiki/Henry_King_(director)
Henry Kissinger	http://en.wikipedia.org/wiki/Henry_Kissinger
Henry Koster	http://en.wikipedia.org/wiki/Henry_Koster
Henry L. Stimson	http://en.wikipedia.org/wiki/Henry_L._Stimson
Henry Laurens	http://en.wikipedia.org/wiki/Henry_Laurens
Henry Laurens Dawes	http://en.wikipedia.org/wiki/Henry_Laurens_Dawes
Henry Lee Lucas	http://en.wikipedia.org/wiki/Henry_Lee_Lucas
Henry Levin	http://en.wikipedia.org/wiki/Henry_Levin
Henry Louis Gates, Jr.	http://en.wikipedia.org/wiki/Henry_Louis_Gates%2C_Jr.
Henry M. Paulson	http://en.wikipedia.org/wiki/Henry_M._Paulson
Henry Mancini	http://en.wikipedia.org/wiki/Henry_Mancini
Henry Mayhew	http://en.wikipedia.org/wiki/Henry_Mayhew
Henry McCullough	http://en.wikipedia.org/wiki/Henry_McCullough
Henry Miller	http://en.wikipedia.org/wiki/Henry_Miller
Henry Moore	http://en.wikipedia.org/wiki/Henry_Moore
Henry Morgenthau, Jr.	http://en.wikipedia.org/wiki/Henry_Morgenthau%2C_Jr.
Henry Morton Stanley	http://en.wikipedia.org/wiki/Henry_Morton_Stanley
Henry of Lausanne	http://en.wikipedia.org/wiki/Henry_of_Lausanne
Henry Pelham	http://en.wikipedia.org/wiki/Henry_Pelham
Henry Petroski	http://en.wikipedia.org/wiki/Henry_Petroski
Henry Purcell	http://en.wikipedia.org/wiki/Henry_Purcell
Henry R. Luce	http://en.wikipedia.org/wiki/Henry_R._Luce
Henry R. Silverman	http://en.wikipedia.org/wiki/Henry_R._Silverman
Henry Richard Vassall Fox	http://en.wikipedia.org/wiki/Henry_Richard_Vassall_Fox
Henry Rollins	http://en.wikipedia.org/wiki/Henry_Rollins
Henry Roth	http://en.wikipedia.org/wiki/Henry_Roth
Henry Sidgwick	http://en.wikipedia.org/wiki/Henry_Sidgwick
Henry Silva	http://en.wikipedia.org/wiki/Henry_Silva
Henry Sloane Coffin	http://en.wikipedia.org/wiki/Henry_Sloane_Coffin
Henry Smith	http://en.wikipedia.org/wiki/Henry_Smith_(British_politician)
Henry Spelman	http://en.wikipedia.org/wiki/Henry_Spelman
Henry Steele Commager	http://en.wikipedia.org/wiki/Henry_Steele_Commager
Henry Stuart Foote	http://en.wikipedia.org/wiki/Henry_Stuart_Foote
Henry Taube	http://en.wikipedia.org/wiki/Henry_Taube
Henry the Navigator	http://en.wikipedia.org/wiki/Henry_the_Navigator
Henry Thomas	http://en.wikipedia.org/wiki/Henry_Thomas
Henry Threadgill	http://en.wikipedia.org/wiki/Henry_Threadgill
Henry van Dyke	http://en.wikipedia.org/wiki/Henry_van_Dyke
Henry Vaughan	http://en.wikipedia.org/wiki/Henry_Vaughan
Henry Vieuxtemps	http://en.wikipedia.org/wiki/Henry_Vieuxtemps
Henry W. Halleck	http://en.wikipedia.org/wiki/Henry_W._Halleck
Henry W. Kendall	http://en.wikipedia.org/wiki/Henry_W._Kendall
Henry Wadsworth Longfellow	http://en.wikipedia.org/wiki/Henry_Wadsworth_Longfellow
Henry Ward Beecher	http://en.wikipedia.org/wiki/Henry_Ward_Beecher
Henry Watterson	http://en.wikipedia.org/wiki/Henry_Watterson
Henry Waxman	http://en.wikipedia.org/wiki/Henry_Waxman
Henry Whitney Bellows	http://en.wikipedia.org/wiki/Henry_Whitney_Bellows
Henry Wilson	http://en.wikipedia.org/wiki/Henry_Wilson
Henry Winkler	http://en.wikipedia.org/wiki/Henry_Winkler
Henry Winter Davis	http://en.wikipedia.org/wiki/Henry_Winter_Davis
Henryk Wieniawski	http://en.wikipedia.org/wiki/Henryk_Wieniawski
Heraclides Ponticus	http://en.wikipedia.org/wiki/Heraclides_Ponticus
Herb Alpert	http://en.wikipedia.org/wiki/Herb_Alpert
Herb Caen	http://en.wikipedia.org/wiki/Herb_Caen
Herb Kelleher	http://en.wikipedia.org/wiki/Herb_Kelleher
Herb Kohl	http://en.wikipedia.org/wiki/Herb_Kohl
Herbert A. Hauptman	http://en.wikipedia.org/wiki/Herbert_A._Hauptman
Herbert A. Simon	http://en.wikipedia.org/wiki/Herbert_A._Simon
Herbert Baxter Adams	http://en.wikipedia.org/wiki/Herbert_Baxter_Adams
Herbert C. Brown	http://en.wikipedia.org/wiki/Herbert_C._Brown
Herbert Fleishhacker	http://en.wikipedia.org/wiki/Herbert_Fleishhacker
Herbert G. Klein	http://en.wikipedia.org/wiki/Herbert_G._Klein
Herbert H. Bateman	http://en.wikipedia.org/wiki/Herbert_H._Bateman
Herbert Henry Asquith	http://en.wikipedia.org/wiki/Herbert_Henry_Asquith
Herbert Hoover	http://en.wikipedia.org/wiki/Herbert_Hoover
Herbert Kroemer	http://en.wikipedia.org/wiki/Herbert_Kroemer
Herbert L. Henkel	http://en.wikipedia.org/wiki/Herbert_L._Henkel
Herbert Lom	http://en.wikipedia.org/wiki/Herbert_Lom
Herbert Marcuse	http://en.wikipedia.org/wiki/Herbert_Marcuse
Herbert Marshall	http://en.wikipedia.org/wiki/Herbert_Marshall
Herbert O. Yardley	http://en.wikipedia.org/wiki/Herbert_O._Yardley
Herbert of Cherbury	http://en.wikipedia.org/wiki/Herbert_of_Cherbury
Herbert Ross	http://en.wikipedia.org/wiki/Herbert_Ross
Herbert S. Zim	http://en.wikipedia.org/wiki/Herbert_S._Zim
Herbert Spencer	http://en.wikipedia.org/wiki/Herbert_Spencer
Herbert Stein	http://en.wikipedia.org/wiki/Herbert_Stein
Herbert Stothart	http://en.wikipedia.org/wiki/Herbert_Stothart
Herbie Hancock	http://en.wikipedia.org/wiki/Herbie_Hancock
Herbie Mann	http://en.wikipedia.org/wiki/Herbie_Mann
Herman Hollerith	http://en.wikipedia.org/wiki/Herman_Hollerith
Herman Melville	http://en.wikipedia.org/wiki/Herman_Melville
Herman Wouk	http://en.wikipedia.org/wiki/Herman_Wouk
Hermann Busenbaum	http://en.wikipedia.org/wiki/Hermann_Busenbaum
Hermann Goering	http://en.wikipedia.org/wiki/Hermann_Goering
Hermann Hesse	http://en.wikipedia.org/wiki/Hermann_Hesse
Hermann Kesten	http://en.wikipedia.org/wiki/Hermann_Kesten
Hermann Mueller	http://en.wikipedia.org/wiki/Hermann_Müller_(politician)
Hermann Nitsch	http://en.wikipedia.org/wiki/Hermann_Nitsch
Hermann Staudinger	http://en.wikipedia.org/wiki/Hermann_Staudinger
Hermann von Helmholtz	http://en.wikipedia.org/wiki/Hermann_von_Helmholtz
Hernando Cortes	http://en.wikipedia.org/wiki/Hernando_Cortes
Hernando de Soto	http://en.wikipedia.org/wiki/Hernando_de_Soto
Hero of Alexandria	http://en.wikipedia.org/wiki/Hero_of_Alexandria
Herod Antipas	http://en.wikipedia.org/wiki/Herod_Antipas
Herod the Great	http://en.wikipedia.org/wiki/Herod_the_Great
Herschel Bernardi	http://en.wikipedia.org/wiki/Herschel_Bernardi
Herschel Walker	http://en.wikipedia.org/wiki/Herschel_Walker
Herschelle Gibbs	http://en.wikipedia.org/wiki/Herschelle_Gibbs
Herv� Villechaize	http://en.wikipedia.org/wiki/Herv%E9_Villechaize
Hervey Allen	http://en.wikipedia.org/wiki/Hervey_Allen
Heston Blumenthal	http://en.wikipedia.org/wiki/Heston_Blumenthal
Hiam Abbass	http://en.wikipedia.org/wiki/Hiam_Abbass
Hideki Saijo	http://en.wikipedia.org/wiki/Hideki_Saijo
Hideki Shirakawa	http://en.wikipedia.org/wiki/Hideki_Shirakawa
Hideki Tojo	http://en.wikipedia.org/wiki/Hideki_Tojo
Hideki Yukawa	http://en.wikipedia.org/wiki/Hideki_Yukawa
Hieronymus Bock	http://en.wikipedia.org/wiki/Hieronymus_Bock
Hieronymus Bosch	http://en.wikipedia.org/wiki/Hieronymus_Bosch
Hifikepunye Pohamba	http://en.wikipedia.org/wiki/Hifikepunye_Pohamba
Hilaire Belloc	http://en.wikipedia.org/wiki/Hilaire_Belloc
Hilarie Burton	http://en.wikipedia.org/wiki/Hilarie_Burton
Hilary Benn	http://en.wikipedia.org/wiki/Hilary_Benn
Hilary Duff	http://en.wikipedia.org/wiki/Hilary_Duff
Hilary Putnam	http://en.wikipedia.org/wiki/Hilary_Putnam
Hilary Rosen	http://en.wikipedia.org/wiki/Hilary_Rosen
Hilary Swank	http://en.wikipedia.org/wiki/Hilary_Swank
Hilda Solis	http://en.wikipedia.org/wiki/Hilda_Solis
Hildegard von Bingen	http://en.wikipedia.org/wiki/Hildegard_von_Bingen
Hill Harper	http://en.wikipedia.org/wiki/Hill_Harper
Hillary Clinton	http://en.wikipedia.org/wiki/Hillary_Clinton
Hillel Slovak	http://en.wikipedia.org/wiki/Hillel_Slovak
Hilmar Orn Hilmarsson	http://en.wikipedia.org/wiki/Hilmar_Orn_Hilmarsson
Hilton Kramer	http://en.wikipedia.org/wiki/Hilton_Kramer
Hines Ward	http://en.wikipedia.org/wiki/Hines_Ward
Hinton Battle	http://en.wikipedia.org/wiki/Hinton_Battle
Hippias of Elis	http://en.wikipedia.org/wiki/Hippias_of_Elis
Hippolyte Taine	http://en.wikipedia.org/wiki/Hippias_of_Elis
Hiram Bingham	http://en.wikipedia.org/wiki/Hiram_Bingham_III
Hiram Fong	http://en.wikipedia.org/wiki/Hiram_Fong
Hiram Johnson	http://en.wikipedia.org/wiki/Hiram_Johnson
Hironari Amano	http://en.wikipedia.org/wiki/Hironari_Amano
Hironobu Sakaguchi	http://en.wikipedia.org/wiki/Hironobu_Sakaguchi
Hiroyuki Sakai	http://en.wikipedia.org/wiki/Hiroyuki_Sakai
Hjalmar Branting	http://en.wikipedia.org/wiki/Hjalmar_Branting
Hjalmar Schacht	http://en.wikipedia.org/wiki/Hjalmar_Schacht
Ho Chi Minh	http://en.wikipedia.org/wiki/Ho_Chi_Minh
Hoagy Carmichael	http://en.wikipedia.org/wiki/Hoagy_Carmichael
Hodding Carter	http://en.wikipedia.org/wiki/Hodding_Carter
Hodding Carter III	http://en.wikipedia.org/wiki/Hodding_Carter_III
Holger Czukay	http://en.wikipedia.org/wiki/Holger_Czukay
Holland Taylor	http://en.wikipedia.org/wiki/Holland_Taylor
Holly Hunter	http://en.wikipedia.org/wiki/Holly_Hunter
Holly Johnson	http://en.wikipedia.org/wiki/Holly_Johnson
Holly Marie Combs	http://en.wikipedia.org/wiki/Holly_Marie_Combs
Holly Robinson Peete	http://en.wikipedia.org/wiki/Holly_Robinson_Peete
Holly Valance	http://en.wikipedia.org/wiki/Holly_Valance
Honor Blackman	http://en.wikipedia.org/wiki/Honor_Blackman
Honor� Daumier	http://en.wikipedia.org/wiki/Honor%E9_Daumier
Honor� de Balzac	http://en.wikipedia.org/wiki/Honor%E9_de_Balzac
Honus Wagner	http://en.wikipedia.org/wiki/Honus_Wagner
Hoot Gibson	http://en.wikipedia.org/wiki/Hoot_Gibson
Hope Davis	http://en.wikipedia.org/wiki/Hope_Davis
Hope Emerson	http://en.wikipedia.org/wiki/Hope_Emerson
Hope Lange	http://en.wikipedia.org/wiki/Hope_Lange
Hope Sandoval	http://en.wikipedia.org/wiki/Hope_Sandoval
Horace Bushnell	http://en.wikipedia.org/wiki/Horace_Bushnell
Horace Greeley	http://en.wikipedia.org/wiki/Horace_Greeley
Horace Gregory	http://en.wikipedia.org/wiki/Horace_Gregory
Horace Liveright	http://en.wikipedia.org/wiki/Horace_Liveright
Horace Mann	http://en.wikipedia.org/wiki/Horace_Mann
Horace Porter	http://en.wikipedia.org/wiki/Horace_Porter
Horace Silver	http://en.wikipedia.org/wiki/Horace_Silver
Horace Walpole	http://en.wikipedia.org/wiki/Horace_Walpole
Horatio Alger	http://en.wikipedia.org/wiki/Horatio_Alger
Horatio Gates	http://en.wikipedia.org/wiki/Horatio_Gates
Horatio Hale	http://en.wikipedia.org/wiki/Horatio_Hale
Horatio Sanz	http://en.wikipedia.org/wiki/Horatio_Sanz
Horst K�hler	http://en.wikipedia.org/wiki/Horst_K%F6hler
Horst K�hler	http://en.wikipedia.org/wiki/Horst_K%F6hler
Horst L. St�rmer	http://en.wikipedia.org/wiki/Horst_L._St%F6rmer
Horst Wessel	http://en.wikipedia.org/wiki/Horst_Wessel
Hortense Calisher	http://en.wikipedia.org/wiki/Hortense_Calisher
Hosni Mubarak	http://en.wikipedia.org/wiki/Hosni_Mubarak
Hosni Mubarak	http://en.wikipedia.org/wiki/Hosni_Mubarak
Hossein Alizadeh	http://en.wikipedia.org/wiki/Hossein_Alizadeh
Hossein Amini	http://en.wikipedia.org/wiki/Hossein_Amini
Howard Ahmanson, Jr.	http://en.wikipedia.org/wiki/Howard_Ahmanson%2C_Jr.
Howard Baker	http://en.wikipedia.org/wiki/Howard_Baker
Howard Berman	http://en.wikipedia.org/wiki/Howard_Berman
Howard Bernstein	http://en.wikipedia.org/wiki/Howard_Bernstein
Howard C. Nielson	http://en.wikipedia.org/wiki/Howard_C._Nielson
Howard Carter	http://en.wikipedia.org/wiki/Howard_Carter
Howard Coble	http://en.wikipedia.org/wiki/Howard_Coble
Howard Coble	http://en.wikipedia.org/wiki/Howard_Coble
Howard Cosell	http://en.wikipedia.org/wiki/Howard_Cosell
Howard Da Silva	http://en.wikipedia.org/wiki/Howard_Da_Silva
Howard Dean	http://en.wikipedia.org/wiki/Howard_Dean
Howard Deutch	http://en.wikipedia.org/wiki/Howard_Deutch
Howard Devoto	http://en.wikipedia.org/wiki/Howard_Devoto
Howard Duff	http://en.wikipedia.org/wiki/Howard_Duff
Howard E. Rollins, Jr.	http://en.wikipedia.org/wiki/Howard_E._Rollins%2C_Jr.
Howard Fast	http://en.wikipedia.org/wiki/Howard_Fast
Howard Fineman	http://en.wikipedia.org/wiki/Howard_Fineman
Howard Hanson	http://en.wikipedia.org/wiki/Howard_Hanson
Howard Hawks	http://en.wikipedia.org/wiki/Howard_Hawks
Howard Hesseman	http://en.wikipedia.org/wiki/Howard_Hesseman
Howard Hughes	http://en.wikipedia.org/wiki/Howard_Hughes
Howard Jarvis	http://en.wikipedia.org/wiki/Howard_Jarvis
Howard Jones	http://en.wikipedia.org/wiki/Howard_Jones_(musician)
Howard K. Smith	http://en.wikipedia.org/wiki/Howard_K._Smith
Howard K. Stern	http://en.wikipedia.org/wiki/Howard_K._Stern
Howard Kaloogian	http://en.wikipedia.org/wiki/Howard_Kaloogian
Howard Keel	http://en.wikipedia.org/wiki/Howard_Keel
Howard Kurtz	http://en.wikipedia.org/wiki/Howard_Kurtz
Howard L. Berman	http://en.wikipedia.org/wiki/Howard_L._Berman
Howard Lindsay	http://en.wikipedia.org/wiki/Howard_Lindsay
Howard Lyman	http://en.wikipedia.org/wiki/Howard_Lyman
Howard M. Metzenbaum	http://en.wikipedia.org/wiki/Howard_M._Metzenbaum
Howard Metzenbaum	http://en.wikipedia.org/wiki/Howard_Metzenbaum
Howard Morris	http://en.wikipedia.org/wiki/Howard_Morris
Howard Moss	http://en.wikipedia.org/wiki/Howard_Moss
Howard Nemerov	http://en.wikipedia.org/wiki/Howard_Nemerov
Howard Pyle	http://en.wikipedia.org/wiki/Howard_Pyle
Howard Rheingold	http://en.wikipedia.org/wiki/Howard_Rheingold
Howard Schultz	http://en.wikipedia.org/wiki/Howard_Schultz
Howard Stern	http://en.wikipedia.org/wiki/Howard_Stern
Howard Sutherland	http://en.wikipedia.org/wiki/Howard_Sutherland
Howard Wolpe	http://en.wikipedia.org/wiki/Howard_Wolpe
Howard Zinn	http://en.wikipedia.org/wiki/Howard_Zinn
Howell Heflin	http://en.wikipedia.org/wiki/Howell_Heflin
Howell Raines	http://en.wikipedia.org/wiki/Howell_Raines
Howell T. Heflin	http://en.wikipedia.org/wiki/Howell_T._Heflin
Howie Carr	http://en.wikipedia.org/wiki/Howie_Carr
Howie D	http://en.wikipedia.org/wiki/Howie_D
Howie Day	http://en.wikipedia.org/wiki/Howie_Day
Howie Long	http://en.wikipedia.org/wiki/Howie_Long
Howie Mandel	http://en.wikipedia.org/wiki/Howie_Mandel
Howlin' Wolf	http://en.wikipedia.org/wiki/Howlin%27_Wolf
Hoyt Axton	http://en.wikipedia.org/wiki/Hoyt_Axton
Hoyt Vandenberg	http://en.wikipedia.org/wiki/Hoyt_Vandenberg
Hoyt Wilhelm	http://en.wikipedia.org/wiki/Hoyt_Wilhelm
Hu Jintao	http://en.wikipedia.org/wiki/Hu_Jintao
Hu Yaobang	http://en.wikipedia.org/wiki/Hu_Yaobang
Hua Guofeng	http://en.wikipedia.org/wiki/Hua_Guofeng
Huang Yong	http://en.wikipedia.org/wiki/Huang_Yong
Hubert de Burgh	http://en.wikipedia.org/wiki/Hubert_de_Burgh
Hubert Howe Bancroft	http://en.wikipedia.org/wiki/Hubert_Howe_Bancroft
Hubert Humphrey	http://en.wikipedia.org/wiki/Hubert_Humphrey
Hubert Ingraham	http://en.wikipedia.org/wiki/Hubert_Ingraham
Hubert Selby	http://en.wikipedia.org/wiki/Hubert_Selby
Hubert Walter	http://en.wikipedia.org/wiki/Hubert_Walter
Huell Howser	http://en.wikipedia.org/wiki/Huell_Howser
Huey Lewis	http://en.wikipedia.org/wiki/Huey_Lewis
Huey Long	http://en.wikipedia.org/wiki/Huey_Long
Huey Newton	http://en.wikipedia.org/wiki/Huey_Newton
Hugh Bayley	http://en.wikipedia.org/wiki/Hugh_Bayley
Hugh Beaumont	http://en.wikipedia.org/wiki/Hugh_Beaumont
Hugh Capet	http://en.wikipedia.org/wiki/Hugh_Capet
Hugh Dancy	http://en.wikipedia.org/wiki/Hugh_Dancy
Hugh Downs	http://en.wikipedia.org/wiki/Hugh_Downs
Hugh Grant	http://en.wikipedia.org/wiki/Hugh_Grant
Hugh Griffith	http://en.wikipedia.org/wiki/Hugh_Griffith
Hugh Hefner	http://en.wikipedia.org/wiki/Hugh_Hefner
Hugh Hopper	http://en.wikipedia.org/wiki/Hugh_Hopper
Hugh Jackman	http://en.wikipedia.org/wiki/Hugh_Jackman
Hugh Kenner	http://en.wikipedia.org/wiki/Hugh_Kenner
Hugh L. Carey	http://en.wikipedia.org/wiki/Hugh_L._Carey
Hugh Latimer	http://en.wikipedia.org/wiki/Hugh_Latimer
Hugh Laurie	http://en.wikipedia.org/wiki/Hugh_Laurie
Hugh le Despenser	http://en.wikipedia.org/wiki/Hugh_Despenser_the_younger
Hugh Lofting	http://en.wikipedia.org/wiki/Hugh_Lofting
Hugh MacDiarmid	http://en.wikipedia.org/wiki/Hugh_MacDiarmid
Hugh MacLennan	http://en.wikipedia.org/wiki/Hugh_MacLennan
Hugh O'Brian	http://en.wikipedia.org/wiki/Hugh_O%27Brian
Hugh O'Neill	http://en.wikipedia.org/wiki/Hugh_O'Neill,_2nd_Earl_of_Tyrone
Hugh Robertson	http://en.wikipedia.org/wiki/Hugh_Robertson_(politician)
Hugh Shelton	http://en.wikipedia.org/wiki/Hugh_Shelton
Hugh Trevor-Roper	http://en.wikipedia.org/wiki/Hugh_Trevor-Roper
Hugo Black	http://en.wikipedia.org/wiki/Hugo_Black
Hugo Chavez	http://en.wikipedia.org/wiki/Hugo_Chavez
Hugo Gernsback	http://en.wikipedia.org/wiki/Hugo_Gernsback
Hugo Grotius	http://en.wikipedia.org/wiki/Hugo_Grotius
Hugo S�nchez	http://en.wikipedia.org/wiki/Hugo_S%E1nchez
Hugo Swire	http://en.wikipedia.org/wiki/Hugo_Swire
Hugo van der Goes	http://en.wikipedia.org/wiki/Hugo_van_der_Goes
Hugo Weaving	http://en.wikipedia.org/wiki/Hugo_Weaving
Hugo Wolf	http://en.wikipedia.org/wiki/Hugo_Wolf
Huldrych Zwingli	http://en.wikipedia.org/wiki/Huldrych_Zwingli
Hulk Hogan	http://en.wikipedia.org/wiki/Hulk_Hogan
Hume Alexander Horan	http://en.wikipedia.org/wiki/Hume_Alexander_Horan
Hume Cronyn	http://en.wikipedia.org/wiki/Hume_Cronyn
Humphrey Bogart	http://en.wikipedia.org/wiki/Humphrey_Bogart
Humphry Davy	http://en.wikipedia.org/wiki/Humphry_Davy
Humphry Osmond	http://en.wikipedia.org/wiki/Humphry_Osmond
Hun Sen	http://en.wikipedia.org/wiki/Hun_Sen
Hunter S. Thompson	http://en.wikipedia.org/wiki/Hunter_S._Thompson
Hunter Tylo	http://en.wikipedia.org/wiki/Hunter_Tylo
Huntz Hall	http://en.wikipedia.org/wiki/Huntz_Hall
Hurricane Carter	http://en.wikipedia.org/wiki/Hurricane_Carter
Husband E. Kimmel	http://en.wikipedia.org/wiki/Husband_E._Kimmel
Hutton Gibson	http://en.wikipedia.org/wiki/Hutton_Gibson
Huw Irranca-Davies	http://en.wikipedia.org/wiki/Huw_Irranca-Davies
Hy Averback	http://en.wikipedia.org/wiki/Hy_Averback
Hyman Rickover	http://en.wikipedia.org/wiki/Hyman_Rickover
Hypatia of Alexandria	http://en.wikipedia.org/wiki/Hypatia_of_Alexandria
Hywel Francis	http://en.wikipedia.org/wiki/Hywel_Francis
Hywel Williams	http://en.wikipedia.org/wiki/Hywel_Williams
I. A. Richards	http://en.wikipedia.org/wiki/I._A._Richards
I. F. Stone	http://en.wikipedia.org/wiki/I._F._Stone
I. M. Pei	http://en.wikipedia.org/wiki/I._M._Pei
Iain Banks	http://en.wikipedia.org/wiki/Iain_Banks
Iain Duncan Smith	http://en.wikipedia.org/wiki/Iain_Duncan_Smith
Iain Sinclair	http://en.wikipedia.org/wiki/Iain_Sinclair
Iain Stewart	http://en.wikipedia.org/wiki/Iain_Stewart_(politician)
Iain Wright	http://en.wikipedia.org/wiki/Iain_Wright
Iajuddin Ahmed	http://en.wikipedia.org/wiki/Iajuddin_Ahmed
Ian Anderson	http://en.wikipedia.org/wiki/Ian_Anderson_(musician)
Ian Austin	http://en.wikipedia.org/wiki/Ian_Austin_(politician)
Ian Bairnson	http://en.wikipedia.org/wiki/Ian_Bairnson
Ian Botham	http://en.wikipedia.org/wiki/Ian_Botham
Ian Brady	http://en.wikipedia.org/wiki/Ian_Brady
Ian Brown	http://en.wikipedia.org/wiki/Ian_Brown
Ian Carmichael	http://en.wikipedia.org/wiki/Ian_Carmichael
Ian Curtis	http://en.wikipedia.org/wiki/Ian_Curtis
Ian Davidson	http://en.wikipedia.org/wiki/Ian_Davidson_(Scottish_politician)
Ian Dury	http://en.wikipedia.org/wiki/Ian_Dury
Ian Fleming	http://en.wikipedia.org/wiki/Ian_Fleming
Ian Gillan	http://en.wikipedia.org/wiki/Ian_Gillan
Ian Hart	http://en.wikipedia.org/wiki/Ian_Hart
Ian Holm	http://en.wikipedia.org/wiki/Ian_Holm
Ian Hunter	http://en.wikipedia.org/wiki/Ian_Hunter_(singer)
Ian Huntley	http://en.wikipedia.org/wiki/Ian_Huntley
Ian Khama	http://en.wikipedia.org/wiki/Ian_Khama
Ian Lavery	http://en.wikipedia.org/wiki/Ian_Lavery
Ian Liddell-Grainger	http://en.wikipedia.org/wiki/Ian_Liddell-Grainger
Ian Lucas	http://en.wikipedia.org/wiki/Ian_Lucas
Ian MacKaye	http://en.wikipedia.org/wiki/Ian_MacKaye
Ian McCulloch	http://en.wikipedia.org/wiki/Ian_McCulloch_(singer)
Ian McDiarmid	http://en.wikipedia.org/wiki/Ian_McDiarmid
Ian McDonald	http://en.wikipedia.org/wiki/Ian_McDonald_(musician)
Ian McEwan	http://en.wikipedia.org/wiki/Ian_McEwan
Ian McKellen	http://en.wikipedia.org/wiki/Ian_McKellen
Ian McLagan	http://en.wikipedia.org/wiki/Ian_McLagan
Ian McShane	http://en.wikipedia.org/wiki/Ian_McShane
Ian Mearns	http://en.wikipedia.org/wiki/Ian_Mearns
Ian Murray	http://en.wikipedia.org/wiki/Ian_Murray_(Scottish_politician)
Ian Paisley Junior	http://en.wikipedia.org/wiki/Ian_Paisley_Junior
Ian Smith	http://en.wikipedia.org/wiki/Ian_Smith
Ian Somerhalder	http://en.wikipedia.org/wiki/Ian_Somerhalder
Ian Swales	http://en.wikipedia.org/wiki/Ian_Swales
Ian Thorpe	http://en.wikipedia.org/wiki/Ian_Thorpe
Ian Underwood	http://en.wikipedia.org/wiki/Ian_Underwood
Ian Wallace	http://en.wikipedia.org/wiki/Ian_Wallace_(drummer)
Ian Wright	http://en.wikipedia.org/wiki/Ian_Wright
Ian Ziering	http://en.wikipedia.org/wiki/Ian_Ziering
Iannis Xenakis	http://en.wikipedia.org/wiki/Iannis_Xenakis
Ibrahim al-Jaafari	http://en.wikipedia.org/wiki/Ibrahim_al-Jaafari
Ibrahim al-Jaafari	http://en.wikipedia.org/wiki/Ibrahim_al-Jaafari
Ibrahim Rugova	http://en.wikipedia.org/wiki/Ibrahim_Rugova
Ibrahim Rugova	http://en.wikipedia.org/wiki/Ibrahim_Rugova
Ice Cube	http://en.wikipedia.org/wiki/Ice_Cube
Iceberg Slim	http://en.wikipedia.org/wiki/Iceberg_Slim
Ida B. Wells-Barnett	http://en.wikipedia.org/wiki/Ida_B._Wells-Barnett
Ida Lupino	http://en.wikipedia.org/wiki/Ida_Lupino
Ida M. Tarbell	http://en.wikipedia.org/wiki/Ida_M._Tarbell
Ida Rentoul Outhwaite	http://en.wikipedia.org/wiki/Ida_Rentoul_Outhwaite
Idi Amin	http://en.wikipedia.org/wiki/Idi_Amin
Idi Amin	http://en.wikipedia.org/wiki/Idi_Amin
Idina Menzel	http://en.wikipedia.org/wiki/Idina_Menzel
Idris Elba	http://en.wikipedia.org/wiki/Idris_Elba
Idriss D�by	http://en.wikipedia.org/wiki/Idriss_D%E9by
Iggy Pop	http://en.wikipedia.org/wiki/Iggy_Pop
Ignace Paderewski	http://en.wikipedia.org/wiki/Ignace_Paderewski
Ignacio Aldecoa	http://en.wikipedia.org/wiki/Ignacio_Aldecoa
Ignacio Milam Tang	http://en.wikipedia.org/wiki/Ignacio_Milam_Tang
Ignatius Donnelly	http://en.wikipedia.org/wiki/Ignatius_Donnelly
Ignatius of Antioch	http://en.wikipedia.org/wiki/Ignatius_of_Antioch
Ignaz Semmelweis	http://en.wikipedia.org/wiki/Ignaz_Semmelweis
Ignazio Silone	http://en.wikipedia.org/wiki/Ignazio_Silone
Igor Ivanov	http://en.wikipedia.org/wiki/Igor_Ivanov
Igor Smirnov	http://en.wikipedia.org/wiki/Igor_Smirnov
Igor Stravinsky	http://en.wikipedia.org/wiki/Igor_Stravinsky
Igor Y. Tamm	http://en.wikipedia.org/wiki/Igor_Y._Tamm
Ike Skelton	http://en.wikipedia.org/wiki/Ike_Skelton
Ike Skelton	http://en.wikipedia.org/wiki/Ike_Skelton
Ike Turner	http://en.wikipedia.org/wiki/Ike_Turner
Ikue Mori	http://en.wikipedia.org/wiki/Ikue_Mori
Ileana Ros-Lehtinen	http://en.wikipedia.org/wiki/Ileana_Ros-Lehtinen
Ilham Aliyev	http://en.wikipedia.org/wiki/Ilham_Aliyev
Ilhan Mimaroglu	http://en.wikipedia.org/wiki/Ilhan_Mimaroglu
Ilie Nastase	http://en.wikipedia.org/wiki/Ilie_Nastase
Illeana Douglas	http://en.wikipedia.org/wiki/Illeana_Douglas
Illinois Jacquet	http://en.wikipedia.org/wiki/Illinois_Jacquet
Ilya Kabakov	http://en.wikipedia.org/wiki/Ilya_Kabakov
Ilya M. Frank	http://en.wikipedia.org/wiki/Ilya_Frank
Ilya Prigogine	http://en.wikipedia.org/wiki/Ilya_Prigogine
Imad Fayez Mugniyah	http://en.wikipedia.org/wiki/Imad_Fayez_Mugniyah
Imelda Marcos	http://en.wikipedia.org/wiki/Imelda_Marcos
Immanuel Kant	http://en.wikipedia.org/wiki/Immanuel_Kant
Immanuel Velikovsky	http://en.wikipedia.org/wiki/Immanuel_Velikovsky
Imogene Coca	http://en.wikipedia.org/wiki/Imogene_Coca
Imran Khan	http://en.wikipedia.org/wiki/Imran_Khan
Imre Kert�sz	http://en.wikipedia.org/wiki/Imre_Kert%E9sz
Imre Nagy	http://en.wikipedia.org/wiki/Imre_Nagy
Increase Mather	http://en.wikipedia.org/wiki/Increase_Mather
Inder Kumar Gujral	http://en.wikipedia.org/wiki/Inder_Kumar_Gujral
India Arie	http://en.wikipedia.org/wiki/India_Arie
Indira Gandhi	http://en.wikipedia.org/wiki/Indira_Gandhi
Inga Swenson	http://en.wikipedia.org/wiki/Inga_Swenson
Inge Meysel	http://en.wikipedia.org/wiki/Inge_Meysel
Inger Stevens	http://en.wikipedia.org/wiki/Inger_Stevens
Ingmar Bergman	http://en.wikipedia.org/wiki/Ingmar_Bergman
Ingrid Bergman	http://en.wikipedia.org/wiki/Ingrid_Bergman
Ingrid Bergman	http://en.wikipedia.org/wiki/Ingrid_Bergman
Ingrid Thulin	http://en.wikipedia.org/wiki/Ingrid_Thulin
Ingvar Kamprad	http://en.wikipedia.org/wiki/Ingvar_Kamprad
Inigo Jones	http://en.wikipedia.org/wiki/Inigo_Jones
Inspecta Deck	http://en.wikipedia.org/wiki/Inspecta_Deck
Inzamam Ul Haq	http://en.wikipedia.org/wiki/Inzamam_Ul_Haq
Ioan Gruffudd	http://en.wikipedia.org/wiki/Ioan_Gruffudd
Iolu Abil	http://en.wikipedia.org/wiki/Iolu_Abil
Ion Aldea-Teodorovici	http://en.wikipedia.org/wiki/Ion_Aldea-Teodorovici
Ion Iliescu	http://en.wikipedia.org/wiki/Ion_Iliescu
Ione Skye	http://en.wikipedia.org/wiki/Ione_Skye
Ira Allen	http://en.wikipedia.org/wiki/Ira_Allen
Ira Einhorn	http://en.wikipedia.org/wiki/Ira_Einhorn
Ira Flatow	http://en.wikipedia.org/wiki/Ira_Flatow
Ira Gershwin	http://en.wikipedia.org/wiki/Ira_Gershwin
Ira Glass	http://en.wikipedia.org/wiki/Ira_Glass
Ira Levin	http://en.wikipedia.org/wiki/Ira_Levin
Ira Magaziner	http://en.wikipedia.org/wiki/Ira_Magaziner
Irene Cara	http://en.wikipedia.org/wiki/Irene_Cara
Irene Dunne	http://en.wikipedia.org/wiki/Irene_Dunne
Ir�ne Joliot-Curie	http://en.wikipedia.org/wiki/Ir%E8ne_Joliot-Curie
Irene Ryan	http://en.wikipedia.org/wiki/Irene_Ryan
Iris Chang	http://en.wikipedia.org/wiki/Iris_Chang
Iris Murdoch	http://en.wikipedia.org/wiki/Iris_Murdoch
Irlene Mandrell	http://en.wikipedia.org/wiki/Irlene_Mandrell
Irma Thomas	http://en.wikipedia.org/wiki/Irma_Thomas
Irv Kupcinet	http://en.wikipedia.org/wiki/Irv_Kupcinet
Irvin Kershner	http://en.wikipedia.org/wiki/Irvin_Kershner
Irvin S. Cobb	http://en.wikipedia.org/wiki/Irvin_S._Cobb
Irvine Welsh	http://en.wikipedia.org/wiki/Irvine_Welsh
Irving Babbitt	http://en.wikipedia.org/wiki/Irving_Babbitt
Irving Berlin	http://en.wikipedia.org/wiki/Irving_Berlin
Irving Fisher	http://en.wikipedia.org/wiki/Irving_Fisher
Irving Howe	http://en.wikipedia.org/wiki/Irving_Howe
Irving Kristol	http://en.wikipedia.org/wiki/Irving_Kristol
Irving Langmuir	http://en.wikipedia.org/wiki/Irving_Langmuir
Irving Mills	http://en.wikipedia.org/wiki/Irving_Mills
Irving Pichel	http://en.wikipedia.org/wiki/Irving_Pichel
Irving Stone	http://en.wikipedia.org/wiki/Irving_Stone
Irving Thalberg	http://en.wikipedia.org/wiki/Irving_Thalberg
Irving Wallace	http://en.wikipedia.org/wiki/Irving_Wallace
Irwin Edman	http://en.wikipedia.org/wiki/Irwin_Edman
Irwin Shaw	http://en.wikipedia.org/wiki/Irwin_Shaw
Isaac Alb�niz	http://en.wikipedia.org/wiki/Isaac_Alb%E9niz
Isaac Asimov	http://en.wikipedia.org/wiki/Isaac_Asimov
Isaac Bashevis Singer	http://en.wikipedia.org/wiki/Isaac_Bashevis_Singer
Isaac ben Solomon Luria	http://en.wikipedia.org/wiki/Isaac_ben_Solomon_Luria
Isaac Brock	http://en.wikipedia.org/wiki/Isaac_Brock_(musician)
Isaac Casaubon	http://en.wikipedia.org/wiki/Isaac_Casaubon
Isaac Chauncey	http://en.wikipedia.org/wiki/Isaac_Chauncey
Isaac da Costa	http://en.wikipedia.org/wiki/Isaac_da_Costa
Isaac Hanson	http://en.wikipedia.org/wiki/Isaac_Hanson
Isaac Hayes	http://en.wikipedia.org/wiki/Isaac_Hayes
Isaac Mizrahi	http://en.wikipedia.org/wiki/Isaac_Mizrahi
Isaac Newton	http://en.wikipedia.org/wiki/Isaac_Newton
Isaac Oliver	http://en.wikipedia.org/wiki/Isaac_Oliver
Isaac Shelby	http://en.wikipedia.org/wiki/Isaac_Shelby
Isaac Stern	http://en.wikipedia.org/wiki/Isaac_Stern
Isabel Allende	http://en.wikipedia.org/wiki/Isabel_Allende
Isabel Peron	http://en.wikipedia.org/wiki/Isabel_Peron
Isabel Sanford	http://en.wikipedia.org/wiki/Isabel_Sanford
Isabella Rossellini	http://en.wikipedia.org/wiki/Isabella_Rossellini
Isabelle Adjani	http://en.wikipedia.org/wiki/Isabelle_Adjani
Isabelle Amyes	http://en.wikipedia.org/wiki/Isabelle_Amyes
Isabelle Huppert	http://en.wikipedia.org/wiki/Isabelle_Huppert
Isadora Duncan	http://en.wikipedia.org/wiki/Isadora_Duncan
Isaiah Berlin	http://en.wikipedia.org/wiki/Isaiah_Berlin
Isaias Afwerki	http://en.wikipedia.org/wiki/Isaias_Afwerki
Ish Kabibble	http://en.wikipedia.org/wiki/Ish_Kabibble
Ishmael Reed	http://en.wikipedia.org/wiki/Ishmael_Reed
Isiah Thomas	http://en.wikipedia.org/wiki/Isiah_Thomas
Isidor Isaac Rabi	http://en.wikipedia.org/wiki/Isidor_Isaac_Rabi
Isidore Mvouba	http://en.wikipedia.org/wiki/Isidore_Mvouba
Isidore of Seville	http://en.wikipedia.org/wiki/Isidore_of_Seville
Isla Blair	http://en.wikipedia.org/wiki/Isla_Blair
Isla Fisher	http://en.wikipedia.org/wiki/Isla_Fisher
Islam Karimov	http://en.wikipedia.org/wiki/Islam_Karimov
Ismail Haniyeh	http://en.wikipedia.org/wiki/Ismail_Haniyeh
Ismail Merchant	http://en.wikipedia.org/wiki/Ismail_Merchant
Ismail Omar Guelleh	http://en.wikipedia.org/wiki/Ismail_Omar_Guelleh
Ismail Pasha	http://en.wikipedia.org/wiki/Ismail_Pasha
Ismet Inonu	http://en.wikipedia.org/wiki/Ismet_Inonu
Isobel Elsom	http://en.wikipedia.org/wiki/Isobel_Elsom
Isoroku Yamamoto	http://en.wikipedia.org/wiki/Isoroku_Yamamoto
Israel Putnam	http://en.wikipedia.org/wiki/Israel_Putnam
Israel Zangwill	http://en.wikipedia.org/wiki/Israel_Zangwill
Isser Harel	http://en.wikipedia.org/wiki/Isser_Harel
Istv�n Sz�chenyi	http://en.wikipedia.org/wiki/Istv%E1n_Sz%E9chenyi
Italo Calvino	http://en.wikipedia.org/wiki/Italo_Calvino
Ito Hirobumi	http://en.wikipedia.org/wiki/Ito_Hirobumi
Itzhak Perlman	http://en.wikipedia.org/wiki/Itzhak_Perlman
Iva Toguri	http://en.wikipedia.org/wiki/Iva_Toguri
Ivan Boesky	http://en.wikipedia.org/wiki/Ivan_Boesky
Ivan Brunetti	http://en.wikipedia.org/wiki/Ivan_Brunetti
Ivan Bunin	http://en.wikipedia.org/wiki/Ivan_Bunin
Ivan G. Seidenberg	http://en.wikipedia.org/wiki/Ivan_G._Seidenberg
Ivan Illich	http://en.wikipedia.org/wiki/Ivan_Illich
Ivan Lendl	http://en.wikipedia.org/wiki/Ivan_Lendl
Ivan Lewis	http://en.wikipedia.org/wiki/Ivan_Lewis
Ivan Pavlov	http://en.wikipedia.org/wiki/Ivan_Pavlov
Ivan Reitman	http://en.wikipedia.org/wiki/Ivan_Reitman
Ivan Rybkin	http://en.wikipedia.org/wiki/Ivan_Rybkin
Ivan Stang	http://en.wikipedia.org/wiki/Ivan_Stang
Ivan the Terrible	http://en.wikipedia.org/wiki/Ivan_the_Terrible
Ivan Turgenev	http://en.wikipedia.org/wiki/Ivan_Turgenev
Ivana Trump	http://en.wikipedia.org/wiki/Ivana_Trump
Ivar Giaever	http://en.wikipedia.org/wiki/Ivar_Giaever
Ivo Sanader	http://en.wikipedia.org/wiki/Ivo_Sanader
Ivo Watts-Russell	http://en.wikipedia.org/wiki/Ivo_Watts-Russell
Ivor Cutler	http://en.wikipedia.org/wiki/Ivor_Cutler
Ivy Compton-Burnett	http://en.wikipedia.org/wiki/Ivy_Compton-Burnett
Ivy Queen	http://en.wikipedia.org/wiki/Ivy_Queen
Iyad Allawi	http://en.wikipedia.org/wiki/Iyad_Allawi
Izaak Walton	http://en.wikipedia.org/wiki/Izaak_Walton
Izzat Ibrahim al-Douri	http://en.wikipedia.org/wiki/Izzat_Ibrahim_al-Douri
Izzy Stradlin	http://en.wikipedia.org/wiki/Izzy_Stradlin
J Dilla	http://en.wikipedia.org/wiki/J_Dilla
J Mascis	http://en.wikipedia.org/wiki/J_Mascis
J. B. Priestley	http://en.wikipedia.org/wiki/J._B._Priestley
J. B. S. Haldane	http://en.wikipedia.org/wiki/J._B._S._Haldane
J. Bennett Johnston	http://en.wikipedia.org/wiki/J._Bennett_Johnston
J. Bennett Johnston	http://en.wikipedia.org/wiki/J._Bennett_Johnston
J. C. Chasez	http://en.wikipedia.org/wiki/J._C._Chasez
J. C. Watts	http://en.wikipedia.org/wiki/J._C._Watts
J. Caleb Boggs	http://en.wikipedia.org/wiki/J._Caleb_Boggs
J. D. Hayworth	http://en.wikipedia.org/wiki/J._D._Hayworth
J. D. Salinger	http://en.wikipedia.org/wiki/J._D._Salinger
J. Danforth Quayle III	http://en.wikipedia.org/wiki/J._Danforth_Quayle_III
J. Edgar Hoover	http://en.wikipedia.org/wiki/J._Edgar_Hoover
J. Franklin Jameson	http://en.wikipedia.org/wiki/J._Franklin_Jameson
J. G. Ballard	http://en.wikipedia.org/wiki/J._G._Ballard
J. G. Thirlwell	http://en.wikipedia.org/wiki/J._G._Thirlwell
J. Georg Bednorz	http://en.wikipedia.org/wiki/J._Georg_Bednorz
J. H. Plumb	http://en.wikipedia.org/wiki/J._H._Plumb
J. Hans D. Jensen	http://en.wikipedia.org/wiki/J._Hans_D._Jensen
J. Hillis Miller	http://en.wikipedia.org/wiki/J._Hillis_Miller
J. I. Packer	http://en.wikipedia.org/wiki/J._I._Packer
J. Irwin Miller	http://en.wikipedia.org/wiki/J._Irwin_Miller
J. J. Cale	http://en.wikipedia.org/wiki/J._J._Cale
J. J. Jackson	http://en.wikipedia.org/wiki/J.J._Jackson_(media_personality)
J. J. Thomson	http://en.wikipedia.org/wiki/J._J._Thomson
J. K. Rowling	http://en.wikipedia.org/wiki/J._K._Rowling
J. K. Simmons	http://en.wikipedia.org/wiki/J._K._Simmons
J. Krishnamurti	http://en.wikipedia.org/wiki/J._Krishnamurti
J. Lee Thompson	http://en.wikipedia.org/wiki/J._Lee_Thompson
J. Leonard Reinsch	http://en.wikipedia.org/wiki/J._Leonard_Reinsch
J. M. Barrie	http://en.wikipedia.org/wiki/J._M._Barrie
J. M. W. Turner	http://en.wikipedia.org/wiki/J._M._W._Turner
J. Otto Seibold	http://en.wikipedia.org/wiki/J._Otto_Seibold
J. P. Donleavy	http://en.wikipedia.org/wiki/J._P._Donleavy
J. Paul Getty, Jr.	http://en.wikipedia.org/wiki/J._Paul_Getty%2C_Jr.
J. Paul Getty, Sr.	http://en.wikipedia.org/wiki/J._Paul_Getty
J. Pierpont Morgan	http://en.wikipedia.org/wiki/J._Pierpont_Morgan
J. R. R. Tolkien	http://en.wikipedia.org/wiki/J._R._R._Tolkien
J. R. Simplot	http://en.wikipedia.org/wiki/J._R._Simplot
J. Roy Rowland	http://en.wikipedia.org/wiki/J._Roy_Rowland
J. T. Money	http://en.wikipedia.org/wiki/JT_Money
J. T. Walsh	http://en.wikipedia.org/wiki/J._T._Walsh
J. Willard Marriott	http://en.wikipedia.org/wiki/J._Willard_Marriott
J. William Fulbright	http://en.wikipedia.org/wiki/J._William_Fulbright
J. Z. Knight	http://en.wikipedia.org/wiki/J._Z._Knight
J.J. Pickle	http://en.wikipedia.org/wiki/J.J._Pickle
Ja Rule	http://en.wikipedia.org/wiki/Ja_Rule
Jaber Al-Ahmad Al-Jaber Al-Sabah	http://en.wikipedia.org/wiki/Jaber_Al-Ahmad_Al-Jaber_Al-Sabah
Jaber III al-Sabah	http://en.wikipedia.org/wiki/Jaber_III_al-Sabah
Jack Abramoff	http://en.wikipedia.org/wiki/Jack_Abramoff
Jack Albertson	http://en.wikipedia.org/wiki/Jack_Albertson
Jack Anderson	http://en.wikipedia.org/wiki/Jack_Anderson_(columnist)
Jack Benny	http://en.wikipedia.org/wiki/Jack_Benny
Jack Black	http://en.wikipedia.org/wiki/Jack_Black
Jack Brooks	http://en.wikipedia.org/wiki/Jack_Brooks_(politician)
Jack Bruce	http://en.wikipedia.org/wiki/Jack_Bruce
Jack Buck	http://en.wikipedia.org/wiki/Jack_Buck
Jack Cafferty	http://en.wikipedia.org/wiki/Jack_Cafferty
Jack Carson	http://en.wikipedia.org/wiki/Jack_Carson
Jack Cassidy	http://en.wikipedia.org/wiki/Jack_Cassidy
Jack Chick	http://en.wikipedia.org/wiki/Jack_Chick
Jack Conway	http://en.wikipedia.org/wiki/Jack_Conway_(filmmaker)
Jack Cope	http://en.wikipedia.org/wiki/Jack_Cope
Jack Dangers	http://en.wikipedia.org/wiki/Jack_Dangers
Jack Davenport	http://en.wikipedia.org/wiki/Jack_Davenport
Jack Dempsey	http://en.wikipedia.org/wiki/Jack_Dempsey
Jack Dromey	http://en.wikipedia.org/wiki/Jack_Dromey
Jack Elam	http://en.wikipedia.org/wiki/Jack_Elam
Jack Fields	http://en.wikipedia.org/wiki/Jack_Fields
Jack Finney	http://en.wikipedia.org/wiki/Jack_Finney
Jack Fletcher	http://en.wikipedia.org/wiki/Jack_Fletcher
Jack Germond	http://en.wikipedia.org/wiki/Jack_Germond
Jack Haley	http://en.wikipedia.org/wiki/Jack_Haley
Jack Hawkins	http://en.wikipedia.org/wiki/Jack_Hawkins
Jack Herer	http://en.wikipedia.org/wiki/Jack_Herer
Jack Holt	http://en.wikipedia.org/wiki/Jack_Holt_(actor)
Jack Idema	http://en.wikipedia.org/wiki/Jack_Idema
Jack Irons	http://en.wikipedia.org/wiki/Jack_Irons
Jack Johnson	http://en.wikipedia.org/wiki/Jack_Johnson_(musician)
Jack Jones	http://en.wikipedia.org/wiki/Jack_Jones_(singer)
Jack Kamen	http://en.wikipedia.org/wiki/Jack_Kamen
Jack Kelley	http://en.wikipedia.org/wiki/Jack_Kelley
Jack Kemp	http://en.wikipedia.org/wiki/Jack_Kemp
Jack Kemp	http://en.wikipedia.org/wiki/Jack_Kemp
Jack Kerouac	http://en.wikipedia.org/wiki/Jack_Kerouac
Jack Kevorkian	http://en.wikipedia.org/wiki/Jack_Kevorkian
Jack Kingston	http://en.wikipedia.org/wiki/Jack_Kingston
Jack Kirby	http://en.wikipedia.org/wiki/Jack_Kirby
Jack Klugman	http://en.wikipedia.org/wiki/Jack_Klugman
Jack L. Chalker	http://en.wikipedia.org/wiki/Jack_L._Chalker
Jack La Lanne	http://en.wikipedia.org/wiki/Jack_La_Lanne
Jack Larson	http://en.wikipedia.org/wiki/Jack_Larson
Jack Lemmon	http://en.wikipedia.org/wiki/Jack_Lemmon
Jack London	http://en.wikipedia.org/wiki/Jack_London
Jack London	http://en.wikipedia.org/wiki/Jack_London
Jack Lopresti	http://en.wikipedia.org/wiki/Jack_Lopresti
Jack Lord	http://en.wikipedia.org/wiki/Jack_Lord
Jack Lynch	http://en.wikipedia.org/wiki/Jack_Lynch
Jack McConnell	http://en.wikipedia.org/wiki/Jack_McConnell
Jack Mullaney	http://en.wikipedia.org/wiki/Jack_Mullaney
Jack Murtha	http://en.wikipedia.org/wiki/Jack_Murtha
Jack Nance	http://en.wikipedia.org/wiki/Jack_Nance
Jack Nicholson	http://en.wikipedia.org/wiki/Jack_Nicholson
Jack Nicklaus	http://en.wikipedia.org/wiki/Jack_Nicklaus
Jack Oakie	http://en.wikipedia.org/wiki/Jack_Oakie
Jack Osbourne	http://en.wikipedia.org/wiki/Jack_Osbourne
Jack Paar	http://en.wikipedia.org/wiki/Jack_Paar
Jack Palance	http://en.wikipedia.org/wiki/Jack_Palance
Jack Parsons	http://en.wikipedia.org/wiki/Jack_Parsons
Jack Quinn	http://en.wikipedia.org/wiki/Jack_Quinn_(politician)
Jack Reed	http://en.wikipedia.org/wiki/Jack_Reed
Jack Roche	http://en.wikipedia.org/wiki/Jack_Roche
Jack Ruby	http://en.wikipedia.org/wiki/Jack_Ruby
Jack S. Kilby	http://en.wikipedia.org/wiki/Jack_S._Kilby
Jack Scalia	http://en.wikipedia.org/wiki/Jack_Scalia
Jack Schmitt	http://en.wikipedia.org/wiki/Jack_Schmitt
Jack Sheppard	http://en.wikipedia.org/wiki/Jack_Sheppard
Jack Soo	http://en.wikipedia.org/wiki/Jack_Soo
Jack Steinberger	http://en.wikipedia.org/wiki/Jack_Steinberger
Jack Straw	http://en.wikipedia.org/wiki/Jack_Straw
Jack Thompson	http://en.wikipedia.org/wiki/Jack_Thompson_(activist)
Jack Valenti	http://en.wikipedia.org/wiki/Jack_Valenti
Jack Vance	http://en.wikipedia.org/wiki/Jack_Vance
Jack W. Buechner	http://en.wikipedia.org/wiki/Jack_Buechner
Jack Wagner	http://en.wikipedia.org/wiki/Jack_Wagner_(actor)
Jack Warden	http://en.wikipedia.org/wiki/Jack_Warden
Jack Watson	http://en.wikipedia.org/wiki/Jack_Watson_(Presidential_adviser)
Jack Webb	http://en.wikipedia.org/wiki/Jack_Webb
Jack Welch	http://en.wikipedia.org/wiki/Jack_Welch
Jack White	http://en.wikipedia.org/wiki/Jack_White_(musician)
Jack Whittaker	http://en.wikipedia.org/wiki/Jack_Whittaker_(lottery_winner)
Jack Wild	http://en.wikipedia.org/wiki/Jack_Wild
Jack Williams	http://en.wikipedia.org/wiki/Jack_Williams_%28American_football%29
Jack�e Harry	http://en.wikipedia.org/wiki/Jack%E9e_Harry
Jackie Chan	http://en.wikipedia.org/wiki/Jackie_Chan
Jackie Collins	http://en.wikipedia.org/wiki/Jackie_Collins
Jackie Coogan	http://en.wikipedia.org/wiki/Jackie_Coogan
Jackie Cooper	http://en.wikipedia.org/wiki/Jackie_Cooper
Jackie DeShannon	http://en.wikipedia.org/wiki/Jackie_DeShannon
Jackie Doyle-Price	http://en.wikipedia.org/wiki/Jackie_Doyle-Price
Jackie Gleason	http://en.wikipedia.org/wiki/Jackie_Gleason
Jackie Jackson	http://en.wikipedia.org/wiki/Jackie_Jackson
Jackie Joyner-Kersee	http://en.wikipedia.org/wiki/Jackie_Joyner-Kersee
Jackie Lane	http://en.wikipedia.org/wiki/Jackie_Lane
Jackie Lomax	http://en.wikipedia.org/wiki/Jackie_Lomax
Jackie Martling	http://en.wikipedia.org/wiki/Jackie_Martling
Jackie Mason	http://en.wikipedia.org/wiki/Jackie_Mason
Jackie Robinson	http://en.wikipedia.org/wiki/Jackie_Robinson
Jackie Speier	http://en.wikipedia.org/wiki/Jackie_Speier
Jackie Stewart	http://en.wikipedia.org/wiki/Jackie_Stewart
Jackie Wilson	http://en.wikipedia.org/wiki/Jackie_Wilson
Jackson Browne	http://en.wikipedia.org/wiki/Jackson_Browne
Jackson Pollock	http://en.wikipedia.org/wiki/Jackson_Pollock
Jaclyn Smith	http://en.wikipedia.org/wiki/Jaclyn_Smith
Jaco Pastorius	http://en.wikipedia.org/wiki/Jaco_Pastorius
Jacob A. Riis	http://en.wikipedia.org/wiki/Jacob_A._Riis
Jacob Abbott	http://en.wikipedia.org/wiki/Jacob_Abbott
Jacob Bigelow	http://en.wikipedia.org/wiki/Jacob_Bigelow
Jacob Epstein	http://en.wikipedia.org/wiki/Jacob_Epstein
Jacob H. Gilbert	http://en.wikipedia.org/wiki/Jacob_H._Gilbert
Jacob Jordaens	http://en.wikipedia.org/wiki/Jacob_Jordaens
Jacob Rees-Mogg	http://en.wikipedia.org/wiki/Jacob_Rees-Mogg
Jacob Zuma	http://en.wikipedia.org/wiki/Jacob_Zuma
Jacobus de Voragine	http://en.wikipedia.org/wiki/Jacobus_de_Voragine
Jacobus H. van 't Hoff	http://en.wikipedia.org/wiki/Jacobus_H._van_%27t_Hoff
Jacoby Shaddix	http://en.wikipedia.org/wiki/Jacoby_Shaddix
Jacopo Della Quercia	http://en.wikipedia.org/wiki/Jacopo_Della_Quercia
Jacopo Palma	http://en.wikipedia.org/wiki/Jacopo_Palma
Jacopo Peri	http://en.wikipedia.org/wiki/Jacopo_Peri
Jacqueline Bisset	http://en.wikipedia.org/wiki/Jacqueline_Bisset
Jacqueline Kennedy Onassis	http://en.wikipedia.org/wiki/Jacqueline_Kennedy_Onassis
Jacqueline McKenzie	http://en.wikipedia.org/wiki/Jacqueline_McKenzie
Jacqueline Susann	http://en.wikipedia.org/wiki/Jacqueline_Susann
Jacques Amand Deslongchamps	http://en.wikipedia.org/wiki/Jacques_Amand_Deslongchamps
Jacques Barzun	http://en.wikipedia.org/wiki/Jacques_Barzun
Jacques Bossuet	http://en.wikipedia.org/wiki/Jacques_Bossuet
Jacques Brel	http://en.wikipedia.org/wiki/Jacques_Brel
Jacques Cartier	http://en.wikipedia.org/wiki/Jacques_Cartier
Jacques Cazotte	http://en.wikipedia.org/wiki/Jacques_Cazotte
Jacques Chirac	http://en.wikipedia.org/wiki/Jacques_Chirac
Jacques Chirac	http://en.wikipedia.org/wiki/Jacques_Chirac
Jacques Cousteau	http://en.wikipedia.org/wiki/Jacques_Cousteau
Jacques d'Amboise	http://en.wikipedia.org/wiki/Jacques_d%27Amboise
Jacques de Larosiere	http://en.wikipedia.org/wiki/Jacques_de_Larosiere
Jacques Delille	http://en.wikipedia.org/wiki/Jacques_Delille
Jacques DeMolay	http://en.wikipedia.org/wiki/Jacques_DeMolay
Jacques Derrida	http://en.wikipedia.org/wiki/Jacques_Derrida
Jacques Dominique Cassini	http://en.wikipedia.org/wiki/Dominique,_comte_de_Cassini
Jacques Dutronc	http://en.wikipedia.org/wiki/Jacques_Dutronc
Jacques Gr�vin	http://en.wikipedia.org/wiki/Jacques_Gr%E9vin
Jacques Ibert	http://en.wikipedia.org/wiki/Jacques_Ibert
Jacques Jasmin	http://en.wikipedia.org/wiki/Jacques_Jasmin
Jacques Kallis	http://en.wikipedia.org/wiki/Jacques_Kallis
Jacques Lacan	http://en.wikipedia.org/wiki/Jacques_Lacan
Jacques Loeb	http://en.wikipedia.org/wiki/Jacques_Loeb
Jacques Maritain	http://en.wikipedia.org/wiki/Jacques_Maritain
Jacques Necker	http://en.wikipedia.org/wiki/Jacques_Necker
Jacques Offenbach	http://en.wikipedia.org/wiki/Jacques_Offenbach
Jacques P�pin	http://en.wikipedia.org/wiki/Jacques_P%E9pin
Jacques Ren� H�bert	http://en.wikipedia.org/wiki/Jacques_Ren%E9_H%E9bert
Jacques Rogge	http://en.wikipedia.org/wiki/Jacques_Rogge
Jacques Sarrazin	http://en.wikipedia.org/wiki/Jacques_Sarrazin
Jacques Sylla	http://en.wikipedia.org/wiki/Jacques_Sylla
Jacques Torres	http://en.wikipedia.org/wiki/Jacques_Torres
Jacques Tourneur	http://en.wikipedia.org/wiki/Jacques_Tourneur
Jacques Verg�s	http://en.wikipedia.org/wiki/Jacques_Verg%E8s
Jacques Villeneuve	http://en.wikipedia.org/wiki/Jacques_Villeneuve
Jacques-Louis David	http://en.wikipedia.org/wiki/Jacques-Louis_David
Jacques-Salomon Hadamard	http://en.wikipedia.org/wiki/Jacques-Salomon_Hadamard
Jada Pinkett Smith	http://en.wikipedia.org/wiki/Jada_Pinkett_Smith
Jade Jagger	http://en.wikipedia.org/wiki/Jade_Jagger
Jadranka Kosor	http://en.wikipedia.org/wiki/Jadranka_Kosor
Jah Wobble	http://en.wikipedia.org/wiki/Jah_Wobble
Jai Rodriguez	http://en.wikipedia.org/wiki/Jai_Rodriguez
Jaime B. Fuster Resident	http://en.wikipedia.org/wiki/Jaime_Fuster
Jaime Cardinal Sin	http://en.wikipedia.org/wiki/Jaime_Cardinal_Sin
Jaime Hernandez	http://en.wikipedia.org/wiki/Jaime_Hernandez
Jaime King	http://en.wikipedia.org/wiki/Jaime_King
Jaime Pressly	http://en.wikipedia.org/wiki/Jaime_Pressly
Jaimee Foxworth	http://en.wikipedia.org/wiki/Jaimee_Foxworth
Jakaya Kikwete	http://en.wikipedia.org/wiki/Jakaya_Kikwete
Jake "The Snake" Roberts	http://en.wikipedia.org/wiki/Jake_%22The_Snake%22_Roberts
Jake Berry	http://en.wikipedia.org/wiki/Jake_Berry
Jake Busey	http://en.wikipedia.org/wiki/Jake_Busey
Jake Epstein	http://en.wikipedia.org/wiki/Jake_Epstein
Jake Garn	http://en.wikipedia.org/wiki/Jake_Garn
Jake Gyllenhaal	http://en.wikipedia.org/wiki/Jake_Gyllenhaal
Jake LaMotta	http://en.wikipedia.org/wiki/Jake_LaMotta
Jake Lloyd	http://en.wikipedia.org/wiki/Jake_Lloyd
Jake Pickle	http://en.wikipedia.org/wiki/Jake_Pickle
Jake Thomas	http://en.wikipedia.org/wiki/Jake_Thomas
Jake Weber	http://en.wikipedia.org/wiki/Jake_Weber
Jakob Boehme	http://en.wikipedia.org/wiki/Jakob_Boehme
Jakob Dylan	http://en.wikipedia.org/wiki/Jakob_Dylan
Jakob Michael Reinhold Lenz	http://en.wikipedia.org/wiki/Jakob_Michael_Reinhold_Lenz
Jalal Talabani	http://en.wikipedia.org/wiki/Jalal_Talabani
Jaleel White	http://en.wikipedia.org/wiki/Jaleel_White
Jam Master Jay	http://en.wikipedia.org/wiki/Jam_Master_Jay
Jamaica Kincaid	http://en.wikipedia.org/wiki/Jamaica_Kincaid
Jamal Abdillah	http://en.wikipedia.org/wiki/Jamal_Abdillah
Jamal Lewis	http://en.wikipedia.org/wiki/Jamal_Lewis
James A. Barcia	http://en.wikipedia.org/wiki/James_A._Barcia
James A. Farley	http://en.wikipedia.org/wiki/James_A._Farley
James A. Herne	http://en.wikipedia.org/wiki/James_A._Herne
James A. Johnson	http://en.wikipedia.org/wiki/James_A._Johnson_(businessman)
James A. Leach	http://en.wikipedia.org/wiki/James_A._Leach
James A. McClure	http://en.wikipedia.org/wiki/James_A._McClure
James A. Michener	http://en.wikipedia.org/wiki/James_A._Michener
James A. Traficant Jr.	http://en.wikipedia.org/wiki/James_A._Traficant_Jr.
James Abdnor	http://en.wikipedia.org/wiki/James_Abdnor
James Acton	http://en.wikipedia.org/wiki/James_Acton
James Agee	http://en.wikipedia.org/wiki/James_Agee
James Alan McPherson	http://en.wikipedia.org/wiki/James_Alan_McPherson
James Aldridge	http://en.wikipedia.org/wiki/James_Aldridge
James Arbuthnot	http://en.wikipedia.org/wiki/James_Arbuthnot
James Arness	http://en.wikipedia.org/wiki/James_Arness
James Avery	http://en.wikipedia.org/wiki/James_Avery_(actor)
James B. Conant	http://en.wikipedia.org/wiki/James_B._Conant
James B. Edwards	http://en.wikipedia.org/wiki/James_B._Edwards
James B. Sumner	http://en.wikipedia.org/wiki/James_B._Sumner
James Baker	http://en.wikipedia.org/wiki/James_Baker
James Baldwin	http://en.wikipedia.org/wiki/James_Baldwin_(writer)
James Bamford	http://en.wikipedia.org/wiki/James_Bamford
James Beard	http://en.wikipedia.org/wiki/James_Beard
James Bernard	http://en.wikipedia.org/wiki/James_Bernard_(composer)
James Best	http://en.wikipedia.org/wiki/James_Best
James Billington	http://en.wikipedia.org/wiki/James_H._Billington
James Blinn	http://en.wikipedia.org/wiki/James_Blinn
James Blish	http://en.wikipedia.org/wiki/James_Blish
James Blunt	http://en.wikipedia.org/wiki/James_Blunt
James Boswell	http://en.wikipedia.org/wiki/James_Boswell
James Bovard	http://en.wikipedia.org/wiki/James_Bovard
James Bowdoin	http://en.wikipedia.org/wiki/James_Bowdoin
James Bradley	http://en.wikipedia.org/wiki/James_Bradley
James Brady	http://en.wikipedia.org/wiki/James_Brady
James Branch Cabell	http://en.wikipedia.org/wiki/James_Branch_Cabell
James Bridges	http://en.wikipedia.org/wiki/James_Bridges
James Brokenshire	http://en.wikipedia.org/wiki/James_Brokenshire
James Brolin	http://en.wikipedia.org/wiki/James_Brolin
James Brown	http://en.wikipedia.org/wiki/James_Brown
James Buchanan	http://en.wikipedia.org/wiki/James_Buchanan
James C. Hagerty	http://en.wikipedia.org/wiki/James_C._Hagerty
James Caan	http://en.wikipedia.org/wiki/James_Caan
James Cagney	http://en.wikipedia.org/wiki/James_Cagney
James Callaghan	http://en.wikipedia.org/wiki/James_Callaghan
James Cameron	http://en.wikipedia.org/wiki/James_Cameron
James Cartwright	http://en.wikipedia.org/wiki/James_Cartwright
James Carville	http://en.wikipedia.org/wiki/James_Carville
James Caviezel	http://en.wikipedia.org/wiki/James_Caviezel
James Chadwick	http://en.wikipedia.org/wiki/James_Chadwick
James Chance	http://en.wikipedia.org/wiki/James_Chance
James Clappison	http://en.wikipedia.org/wiki/James_Clappison
James Clarence Mangan	http://en.wikipedia.org/wiki/James_Clarence_Mangan
James Clavell	http://en.wikipedia.org/wiki/James_Clavell
James Clerk Maxwell	http://en.wikipedia.org/wiki/James_Clerk_Maxwell
James Coburn	http://en.wikipedia.org/wiki/James_Coburn
James Coco	http://en.wikipedia.org/wiki/James_Coco
James Comey	http://en.wikipedia.org/wiki/James_Comey
James Conway	http://en.wikipedia.org/wiki/James_T._Conway
James Cook	http://en.wikipedia.org/wiki/James_Cook
James Crichton	http://en.wikipedia.org/wiki/James_Crichton
James Cromwell	http://en.wikipedia.org/wiki/James_Cromwell
James D. Hodgson	http://en.wikipedia.org/wiki/James_D._Hodgson
James Daly	http://en.wikipedia.org/wiki/James_Daly_(actor)
James D'Arcy	http://en.wikipedia.org/wiki/James_D%27Arcy
James Darren	http://en.wikipedia.org/wiki/James_Darren
James Dean	http://en.wikipedia.org/wiki/James_Dean
James DeBarge	http://en.wikipedia.org/wiki/James_DeBarge
James Denton	http://en.wikipedia.org/wiki/James_Denton
James Dewar	http://en.wikipedia.org/wiki/James_Dewar
James Dickey	http://en.wikipedia.org/wiki/James_Dickey
James Dimon	http://en.wikipedia.org/wiki/James_Dimon
James Dobson	http://en.wikipedia.org/wiki/James_Dobson
James Donald	http://en.wikipedia.org/wiki/James_Donald
James Doohan	http://en.wikipedia.org/wiki/James_Doohan
James Doolittle	http://en.wikipedia.org/wiki/Jimmy_Doolittle
James Douglas	http://en.wikipedia.org/wiki/Jim_Douglas
James Drury	http://en.wikipedia.org/wiki/James_Drury
James Duddridge	http://en.wikipedia.org/wiki/James_Duddridge
James Dunn	http://en.wikipedia.org/wiki/James_Dunn_(actor)
James Dwight Dana	http://en.wikipedia.org/wiki/James_Dwight_Dana
James Dyson	http://en.wikipedia.org/wiki/James_Dyson
James E. Cayne	http://en.wikipedia.org/wiki/James_E._Cayne
James E. Rohr	http://en.wikipedia.org/wiki/Jim_Rohr
James E. Watson	http://en.wikipedia.org/wiki/James_E._Watson
James E. West	http://en.wikipedia.org/wiki/James_E._West_(politician)
James Earl Jones	http://en.wikipedia.org/wiki/James_Earl_Jones
James Earl Ray	http://en.wikipedia.org/wiki/James_Earl_Ray
James Edward Meade	http://en.wikipedia.org/wiki/James_Edward_Meade
James Edward Oglethorpe	http://en.wikipedia.org/wiki/James_Edward_Oglethorpe
James Ellroy	http://en.wikipedia.org/wiki/James_Ellroy
James Ensor	http://en.wikipedia.org/wiki/James_Ensor
James F. Byrnes	http://en.wikipedia.org/wiki/James_F._Byrnes
James Fallows	http://en.wikipedia.org/wiki/James_Fallows
James Farentino	http://en.wikipedia.org/wiki/James_Farentino
James Farmer	http://en.wikipedia.org/wiki/James_L._Farmer,_Jr.
James Fenimore Cooper	http://en.wikipedia.org/wiki/James_Fenimore_Cooper
James Florio	http://en.wikipedia.org/wiki/James_Florio
James Ford Rhodes	http://en.wikipedia.org/wiki/James_Ford_Rhodes
James Fox	http://en.wikipedia.org/wiki/James_Fox
James Franciscus	http://en.wikipedia.org/wiki/James_Franciscus
James Franck	http://en.wikipedia.org/wiki/James_Franck
James Franco	http://en.wikipedia.org/wiki/James_Franco
James Freeman Clarke	http://en.wikipedia.org/wiki/James_Freeman_Clarke
James Frey	http://en.wikipedia.org/wiki/James_Frey
James G. Birney	http://en.wikipedia.org/wiki/James_G._Birney
James G. Blaine	http://en.wikipedia.org/wiki/James_G._Blaine
James Gadsden	http://en.wikipedia.org/wiki/James_Gadsden
James Gammon	http://en.wikipedia.org/wiki/James_Gammon
James Gandolfini	http://en.wikipedia.org/wiki/James_Gandolfini
James Garfield	http://en.wikipedia.org/wiki/James_Garfield
James Garner	http://en.wikipedia.org/wiki/James_Garner
James Gillray	http://en.wikipedia.org/wiki/James_Gillray
James Gould Cozzens	http://en.wikipedia.org/wiki/James_Gould_Cozzens
James Grauerholz	http://en.wikipedia.org/wiki/James_Grauerholz
James Gray	http://en.wikipedia.org/wiki/James_Gray_(politician)
James Gray	http://en.wikipedia.org/wiki/James_Gray_%28politician%29
James Greenwood	http://en.wikipedia.org/wiki/James_C._Greenwood
James Gregory	http://en.wikipedia.org/wiki/James_Gregory_(actor)
James H. Quillen	http://en.wikipedia.org/wiki/James_H._Quillen
James H. Scheuer	http://en.wikipedia.org/wiki/James_H._Scheuer
James H. Scheuer	http://en.wikipedia.org/wiki/James_H._Scheuer
James H. Webb	http://en.wikipedia.org/wiki/James_H._Webb
James Hadley Chase	http://en.wikipedia.org/wiki/James_Hadley_Chase
James Hampton	http://en.wikipedia.org/wiki/James_Hampton_(actor)
James Harlan	http://en.wikipedia.org/wiki/James_Harlan_(senator)
James Harrington	http://en.wikipedia.org/wiki/James_Harrington_(author)
James Harvey Robinson	http://en.wikipedia.org/wiki/James_Harvey_Robinson
James Henry Lane	http://en.wikipedia.org/wiki/James_H._Lane_(politician)
James Herriot	http://en.wikipedia.org/wiki/James_Herriot
James Hetfield	http://en.wikipedia.org/wiki/James_Hetfield
James Hewitt	http://en.wikipedia.org/wiki/James_Hewitt
James Hogg	http://en.wikipedia.org/wiki/James_Hogg
James Hong	http://en.wikipedia.org/wiki/James_Hong
James Horner	http://en.wikipedia.org/wiki/James_Horner
James Hutton	http://en.wikipedia.org/wiki/James_Hutton
James I	http://en.wikipedia.org/wiki/James_I_of_Aragon
James I	http://en.wikipedia.org/wiki/James_I_of_Scotland
James Iha	http://en.wikipedia.org/wiki/James_Iha
James II	http://en.wikipedia.org/wiki/James_II_of_Scotland
James III	http://en.wikipedia.org/wiki/James_III_of_Scotland
James Inhofe	http://en.wikipedia.org/wiki/James_Inhofe
James IV	http://en.wikipedia.org/wiki/James_IV
James Ivory	http://en.wikipedia.org/wiki/James_Ivory_(director)
James J. Florio	http://en.wikipedia.org/wiki/James_J._Florio
James J. Howard	http://en.wikipedia.org/wiki/James_J._Howard
James J. Kilpatrick	http://en.wikipedia.org/wiki/James_J._Kilpatrick
James Jones	http://en.wikipedia.org/wiki/James_Jones_(author)
James Joseph Sylvester	http://en.wikipedia.org/wiki/James_Joseph_Sylvester
James Joyce	http://en.wikipedia.org/wiki/James_Joyce
James K. Hahn	http://en.wikipedia.org/wiki/James_K._Hahn
James Kimsey	http://en.wikipedia.org/wiki/James_Kimsey
James Kirby	http://en.wikipedia.org/wiki/James_Kirby
James Kirkwood	http://en.wikipedia.org/wiki/James_Kirkwood,_Jr.
James Knox Polk	http://en.wikipedia.org/wiki/James_Knox_Polk
James L. Brooks	http://en.wikipedia.org/wiki/James_L._Brooks
James L. Buckley	http://en.wikipedia.org/wiki/James_L._Buckley
James L. Jones	http://en.wikipedia.org/wiki/James_L._Jones
James L. McConaughy	http://en.wikipedia.org/wiki/James_L._McConaughy
James L. Oberstar	http://en.wikipedia.org/wiki/James_L._Oberstar
James Lafferty	http://en.wikipedia.org/wiki/James_Lafferty
James Laughlin	http://en.wikipedia.org/wiki/James_Laughlin
James Lavelle	http://en.wikipedia.org/wiki/James_Lavelle
James Lee Witt	http://en.wikipedia.org/wiki/James_Lee_Witt
James Levine	http://en.wikipedia.org/wiki/James_Levine
James Lipton	http://en.wikipedia.org/wiki/James_Lipton
James Longstreet	http://en.wikipedia.org/wiki/James_Longstreet
James Lovelock	http://en.wikipedia.org/wiki/James_Lovelock
James M. Buchanan	http://en.wikipedia.org/wiki/James_M._Buchanan
James M. Cain	http://en.wikipedia.org/wiki/James_M._Cain
James M. Jeffords	http://en.wikipedia.org/wiki/James_M._Jeffords
James M. Kilts	http://en.wikipedia.org/wiki/James_M._Kilts
James MacArthur	http://en.wikipedia.org/wiki/James_MacArthur
James Mackay	http://en.wikipedia.org/wiki/James_A._Mackay
James Macpherson	http://en.wikipedia.org/wiki/James_Macpherson
James Madison	http://en.wikipedia.org/wiki/James_Madison
James Mangold	http://en.wikipedia.org/wiki/James_Mangold
James Marsden	http://en.wikipedia.org/wiki/James_Marsden
James Marsters	http://en.wikipedia.org/wiki/James_Marsters
James Mason	http://en.wikipedia.org/wiki/James_Mason
James McClatchy	http://en.wikipedia.org/wiki/James_B._McClatchy
James McClure	http://en.wikipedia.org/wiki/James_H._McClure
James McDermott	http://en.wikipedia.org/wiki/Jim_McDermott
James McGovern	http://en.wikipedia.org/wiki/Jim_McGovern
James McGreevey	http://en.wikipedia.org/wiki/James_McGreevey
James McNerney	http://en.wikipedia.org/wiki/James_McNerney
James Merrill	http://en.wikipedia.org/wiki/James_Merrill
James Michel	http://en.wikipedia.org/wiki/James_Michel
James Mill	http://en.wikipedia.org/wiki/James_Mill
James Monroe	http://en.wikipedia.org/wiki/James_Monroe
James Morris	http://en.wikipedia.org/wiki/James_Morris_(British_politician)
James Naughton	http://en.wikipedia.org/wiki/James_Naughton
James O. Richardson	http://en.wikipedia.org/wiki/James_O._Richardson
James Oberstar	http://en.wikipedia.org/wiki/James_Oberstar
James Otis	http://en.wikipedia.org/wiki/James_Otis,_Jr.
James P. Hoffa	http://en.wikipedia.org/wiki/James_P._Hoffa
James P. Mitchell	http://en.wikipedia.org/wiki/James_P._Mitchell
James Paice	http://en.wikipedia.org/wiki/James_Paice
James Parkinson	http://en.wikipedia.org/wiki/James_Parkinson
James Parton	http://en.wikipedia.org/wiki/James_Parton
James Patterson	http://en.wikipedia.org/wiki/James_Patterson
James Prescott Joule	http://en.wikipedia.org/wiki/James_Prescott_Joule
James Purdy	http://en.wikipedia.org/wiki/James_Purdy
James Purefoy	http://en.wikipedia.org/wiki/James_Purefoy
James Quello	http://en.wikipedia.org/wiki/James_Quello
James R. Bath	http://en.wikipedia.org/wiki/James_R._Bath
James R. Jones	http://en.wikipedia.org/wiki/James_R._Jones
James R. Schlesinger	http://en.wikipedia.org/wiki/James_R._Schlesinger
James R. Thompson	http://en.wikipedia.org/wiki/James_R._Thompson
James Rainwater	http://en.wikipedia.org/wiki/James_Rainwater
James Ramsay, Marquess of Dalhousie	http://en.wikipedia.org/wiki/James_Broun-Ramsay,_1st_Marquess_of_Dalhousie
James Randi	http://en.wikipedia.org/wiki/James_Randi
James Redfield	http://en.wikipedia.org/wiki/James_Redfield
James Remar	http://en.wikipedia.org/wiki/James_Remar
James Risen	http://en.wikipedia.org/wiki/James_Risen
James Robertson	http://en.wikipedia.org/wiki/James_Robertson_(judge)
James Robison	http://en.wikipedia.org/wiki/James_Robison
James Rolph, Jr.	http://en.wikipedia.org/wiki/James_Rolph%2C_Jr.
James Russell Lowell	http://en.wikipedia.org/wiki/James_Russell_Lowell
James S. Coleman	http://en.wikipedia.org/wiki/James_Samuel_Coleman
James S. Sherman	http://en.wikipedia.org/wiki/James_S._Sherman
James Sanborn	http://en.wikipedia.org/wiki/James_Sanborn
James Schuyler	http://en.wikipedia.org/wiki/James_Schuyler
James Sharp	http://en.wikipedia.org/wiki/James_E._Sharp
James Sheakley	http://en.wikipedia.org/wiki/James_Sheakley
James Shirley	http://en.wikipedia.org/wiki/James_Shirley
James Sinegal	http://en.wikipedia.org/wiki/James_Sinegal
James Smithson	http://en.wikipedia.org/wiki/James_Smithson
James Spader	http://en.wikipedia.org/wiki/James_Spader
James Stacy	http://en.wikipedia.org/wiki/James_Stacy
James Stewart	http://en.wikipedia.org/wiki/James_Stewart
James Stirling	http://en.wikipedia.org/wiki/James_Stirling_(architect)
James Stirling	http://en.wikipedia.org/wiki/James_Stirling_(mathematician)
James Stockdale	http://en.wikipedia.org/wiki/James_Stockdale
James Syme	http://en.wikipedia.org/wiki/James_Syme
James Symington	http://en.wikipedia.org/wiki/James_W._Symington
James T. Broyhill	http://en.wikipedia.org/wiki/James_T._Broyhill
James T. Farrell	http://en.wikipedia.org/wiki/James_T._Farrell
James Tate	http://en.wikipedia.org/wiki/James_Tate_(writer)
James Taylor	http://en.wikipedia.org/wiki/James_Taylor
James Tenney	http://en.wikipedia.org/wiki/James_Tenney
James Thomas Fields	http://en.wikipedia.org/wiki/James_Thomas_Fields
James Thurber	http://en.wikipedia.org/wiki/James_Thurber
James Tobin	http://en.wikipedia.org/wiki/James_Tobin
James Traficant	http://en.wikipedia.org/wiki/James_Traficant
James Truslow Adams	http://en.wikipedia.org/wiki/James_Truslow_Adams
James Ussher	http://en.wikipedia.org/wiki/James_Ussher
James V	http://en.wikipedia.org/wiki/James_V
James V. Forrestal	http://en.wikipedia.org/wiki/James_V._Forrestal
James V. Hansen	http://en.wikipedia.org/wiki/James_V._Hansen
James Van Allen	http://en.wikipedia.org/wiki/James_Van_Allen
James Van Der Beek	http://en.wikipedia.org/wiki/James_Van_Der_Beek
James Van Praagh	http://en.wikipedia.org/wiki/James_Van_Praagh
James W. Cronin	http://en.wikipedia.org/wiki/James_W._Cronin
James W. McCord, Jr.	http://en.wikipedia.org/wiki/James_W._McCord%2C_Jr.
James W. Owens	http://en.wikipedia.org/wiki/James_W._Owens
James W. Wadsworth, Jr.	http://en.wikipedia.org/wiki/James_W._Wadsworth%2C_Jr.
James Watkins	http://en.wikipedia.org/wiki/James_D._Watkins
James Watson	http://en.wikipedia.org/wiki/James_D._Watson
James Watt	http://en.wikipedia.org/wiki/James_Watt
James Watt	http://en.wikipedia.org/wiki/James_Watt
James Weaver	http://en.wikipedia.org/wiki/Jim_Weaver_(Oregon_politician)
James Weldon Johnson	http://en.wikipedia.org/wiki/James_Weldon_Johnson
James Whale	http://en.wikipedia.org/wiki/James_Whale
James Wharton	http://en.wikipedia.org/wiki/James_Wharton_(UK_politician)
James Whistler	http://en.wikipedia.org/wiki/James_Abbott_McNeill_Whistler
James Whitcomb Riley	http://en.wikipedia.org/wiki/James_Whitcomb_Riley
James Whitmore	http://en.wikipedia.org/wiki/James_Whitmore
James Wilkinson	http://en.wikipedia.org/wiki/James_Wilkinson
James Wilson	http://en.wikipedia.org/wiki/James_Wilson
James Wolcott	http://en.wikipedia.org/wiki/James_Wolcott
James Wolfe	http://en.wikipedia.org/wiki/James_Wolfe
James Wolfensohn	http://en.wikipedia.org/wiki/James_Wolfensohn
James Woods	http://en.wikipedia.org/wiki/James_Woods
James Woolsey	http://en.wikipedia.org/wiki/James_Woolsey
James Worthy	http://en.wikipedia.org/wiki/James_Worthy
James Wright	http://en.wikipedia.org/wiki/James_Wright_(poet)
James. A. McClure	http://en.wikipedia.org/wiki/James_A._McClure
Jameson Parker	http://en.wikipedia.org/wiki/Jameson_Parker
Jameson Thomas	http://en.wikipedia.org/wiki/Jameson_Thomas
Jamey Sheridan	http://en.wikipedia.org/wiki/Jamey_Sheridan
Jami Gertz	http://en.wikipedia.org/wiki/Jami_Gertz
Jamie Bell	http://en.wikipedia.org/wiki/Jamie_Bell
Jamie Farr	http://en.wikipedia.org/wiki/Jamie_Farr
Jamie Foxx	http://en.wikipedia.org/wiki/Jamie_Foxx
Jamie Hyneman	http://en.wikipedia.org/wiki/Jamie_Hyneman
Jamie Kennedy	http://en.wikipedia.org/wiki/Jamie_Kennedy
Jamie L. Whitten	http://en.wikipedia.org/wiki/Jamie_L._Whitten
Jamie Lee Curtis	http://en.wikipedia.org/wiki/Jamie_Lee_Curtis
Jamie Lidell	http://en.wikipedia.org/wiki/Jamie_Lidell
Jamie Lynn Spears	http://en.wikipedia.org/wiki/Jamie_Lynn_Spears
Jamie Muir	http://en.wikipedia.org/wiki/Jamie_Muir
Jamie Oliver	http://en.wikipedia.org/wiki/Jamie_Oliver
Jamie Reed	http://en.wikipedia.org/wiki/Jamie_Reed
Jamie S. Gorelick	http://en.wikipedia.org/wiki/Jamie_S._Gorelick
Jamie Thomas	http://en.wikipedia.org/wiki/Jamie_Thomas
Jamie White	http://en.wikipedia.org/wiki/Jamie_White
Jamie Zawinski	http://en.wikipedia.org/wiki/Jamie_Zawinski
Jamie-Lynn DiScala	http://en.wikipedia.org/wiki/Jamie-Lynn_DiScala
Jan Baptist van Helmont	http://en.wikipedia.org/wiki/Jan_Baptist_van_Helmont
Jan Berry	http://en.wikipedia.org/wiki/Jan_Berry
Jan Crawford Greenburg	http://en.wikipedia.org/wiki/Jan_Crawford_Greenburg
Jan Davidsz de Heem	http://en.wikipedia.org/wiki/Jan_Davidsz_de_Heem
Jan de Bont	http://en.wikipedia.org/wiki/Jan_de_Bont
Jan Egeland	http://en.wikipedia.org/wiki/Jan_Egeland
Jan Fischer	http://en.wikipedia.org/wiki/Jan_Fischer_(politician)
Jan Hammer	http://en.wikipedia.org/wiki/Jan_Hammer
Jan Hendrik Oort	http://en.wikipedia.org/wiki/Jan_Hendrik_Oort
Jan Hooks	http://en.wikipedia.org/wiki/Jan_Hooks
Jan Hus	http://en.wikipedia.org/wiki/Jan_Hus
Jan Josephs van Goyen	http://en.wikipedia.org/wiki/Jan_Josephs_van_Goyen
Jan Mabuse	http://en.wikipedia.org/wiki/Jan_Mabuse
Jan Masaryk	http://en.wikipedia.org/wiki/Jan_Masaryk
Jan Meyers	http://en.wikipedia.org/wiki/Jan_Meyers
Jan Miense Molenaer	http://en.wikipedia.org/wiki/Jan_Miense_Molenaer
Jan Miner	http://en.wikipedia.org/wiki/Jan_Miner
Jan Morris	http://en.wikipedia.org/wiki/Jan_Morris
Jan Peter Balkenende	http://en.wikipedia.org/wiki/Jan_Peter_Balkenende
Jan Schakowsky	http://en.wikipedia.org/wiki/Jan_Schakowsky
Jan Simonsen	http://en.wikipedia.org/wiki/Jan_Simonsen
Jan Smithers	http://en.wikipedia.org/wiki/Jan_Smithers
Jan Smuts	http://en.wikipedia.org/wiki/Jan_Smuts
Jan Steen	http://en.wikipedia.org/wiki/Jan_Steen
Jan Sterling	http://en.wikipedia.org/wiki/Jan_Sterling
Jan Swammerdam	http://en.wikipedia.org/wiki/Jan_Swammerdam
Jan Tarnowski	http://en.wikipedia.org/wiki/Jan_Tarnowski
Jan Tinbergen	http://en.wikipedia.org/wiki/Jan_Tinbergen
Jan van Eyck	http://en.wikipedia.org/wiki/Jan_van_Eyck
Jan Vermeer	http://en.wikipedia.org/wiki/Jan_Vermeer
Jane Addams	http://en.wikipedia.org/wiki/Jane_Addams
Jane Alexander	http://en.wikipedia.org/wiki/Jane_Alexander
Jane Asher	http://en.wikipedia.org/wiki/Jane_Asher
Jane Austen	http://en.wikipedia.org/wiki/Jane_Austen
Jane Badler	http://en.wikipedia.org/wiki/Jane_Badler
Jane Birkin	http://en.wikipedia.org/wiki/Jane_Birkin
Jane Bowles	http://en.wikipedia.org/wiki/Jane_Bowles
Jane Bryant Quinn	http://en.wikipedia.org/wiki/Jane_Bryant_Quinn
Jane Campion	http://en.wikipedia.org/wiki/Jane_Campion
Jane Clayson	http://en.wikipedia.org/wiki/Jane_Clayson
Jane Curtin	http://en.wikipedia.org/wiki/Jane_Curtin
Jane Darwell	http://en.wikipedia.org/wiki/Jane_Darwell
Jane Dee Hull	http://en.wikipedia.org/wiki/Jane_Dee_Hull
Jane Ellison	http://en.wikipedia.org/wiki/Jane_Ellison
Jane Fonda	http://en.wikipedia.org/wiki/Jane_Fonda
Jane Goodall	http://en.wikipedia.org/wiki/Jane_Goodall
Jane Greer	http://en.wikipedia.org/wiki/Jane_Greer
Jane Hall	http://en.wikipedia.org/wiki/Jane_Hall_(journalist)
Jane Harman	http://en.wikipedia.org/wiki/Jane_Harman
Jane Horrocks	http://en.wikipedia.org/wiki/Jane_Horrocks
Jane Kaczmarek	http://en.wikipedia.org/wiki/Jane_Kaczmarek
Jane Krakowski	http://en.wikipedia.org/wiki/Jane_Krakowski
Jane Leeves	http://en.wikipedia.org/wiki/Jane_Leeves
Jane Lynch	http://en.wikipedia.org/wiki/Jane_Lynch
Jane March	http://en.wikipedia.org/wiki/Jane_March
Jane Pauley	http://en.wikipedia.org/wiki/Jane_Pauley
Jane Powell	http://en.wikipedia.org/wiki/Jane_Powell
Jane Rule	http://en.wikipedia.org/wiki/Jane_Rule
Jane Russell	http://en.wikipedia.org/wiki/Jane_Russell
Jane Seymour	http://en.wikipedia.org/wiki/Jane_Seymour_(actress)
Jane Smiley	http://en.wikipedia.org/wiki/Jane_Smiley
Jane Velez-Mitchell	http://en.wikipedia.org/wiki/Jane_Velez-Mitchell
Jane Wiedlin	http://en.wikipedia.org/wiki/Jane_Wiedlin
Jane Withers	http://en.wikipedia.org/wiki/Jane_Withers
Jane Wyatt	http://en.wikipedia.org/wiki/Jane_Wyatt
Jane Wyman	http://en.wikipedia.org/wiki/Jane_Wyman
Janeane Garofalo	http://en.wikipedia.org/wiki/Janeane_Garofalo
Janet Cooke	http://en.wikipedia.org/wiki/Janet_Cooke
Janet Fielding	http://en.wikipedia.org/wiki/Janet_Fielding
Janet Flanner	http://en.wikipedia.org/wiki/Janet_Flanner
Janet Frame	http://en.wikipedia.org/wiki/Janet_Frame
Janet Gaynor	http://en.wikipedia.org/wiki/Janet_Gaynor
Janet Jackson	http://en.wikipedia.org/wiki/Janet_Jackson
Janet Jones	http://en.wikipedia.org/wiki/Janet_Jones
Janet Langhart	http://en.wikipedia.org/wiki/Janet_Langhart
Janet Leigh	http://en.wikipedia.org/wiki/Janet_Leigh
Janet Margolin	http://en.wikipedia.org/wiki/Janet_Margolin
Janet Maslin	http://en.wikipedia.org/wiki/Janet_Maslin
Janet Napolitano	http://en.wikipedia.org/wiki/Janet_Napolitano
Janet Reno	http://en.wikipedia.org/wiki/Janet_Reno
Janet Steiger	http://en.wikipedia.org/wiki/Janet_Steiger
Janet Suzman	http://en.wikipedia.org/wiki/Janet_Suzman
Janette Scott	http://en.wikipedia.org/wiki/Janette_Scott
Jani Lane	http://en.wikipedia.org/wiki/Jani_Lane
Janice Dickinson	http://en.wikipedia.org/wiki/Janice_Dickinson
Janine Turner	http://en.wikipedia.org/wiki/Janine_Turner
Janis Ian	http://en.wikipedia.org/wiki/Janis_Ian
Janis Joplin	http://en.wikipedia.org/wiki/Janis_Joplin
Janis Karpinski	http://en.wikipedia.org/wiki/Janis_Karpinski
Jan-Michael Vincent	http://en.wikipedia.org/wiki/Jan-Michael_Vincent
Jann Wenner	http://en.wikipedia.org/wiki/Jann_Wenner
January Jones	http://en.wikipedia.org/wiki/January_Jones
Jared Fogle	http://en.wikipedia.org/wiki/Jared_Fogle
Jared Leto	http://en.wikipedia.org/wiki/Jared_Leto
Jared Padalecki	http://en.wikipedia.org/wiki/Jared_Padalecki
Jared Polis	http://en.wikipedia.org/wiki/Jared_Polis
Jared Sparks	http://en.wikipedia.org/wiki/Jared_Sparks
Jarl Alfredius	http://en.wikipedia.org/wiki/Jarl_Alfredius
Jaromil Jires	http://en.wikipedia.org/wiki/Jaromil_Jires
Jaron Lanier	http://en.wikipedia.org/wiki/Jaron_Lanier
Jaroslav Hasek	http://en.wikipedia.org/wiki/Jaroslav_Hasek
Jaroslav Heyrovsky	http://en.wikipedia.org/wiki/Jaroslav_Heyrovsky
Jaroslav Seifert	http://en.wikipedia.org/wiki/Jaroslav_Seifert
Jarvis Cocker	http://en.wikipedia.org/wiki/Jarvis_Cocker
Jascha Heifetz	http://en.wikipedia.org/wiki/Jascha_Heifetz
Jasmine Guy	http://en.wikipedia.org/wiki/Jasmine_Guy
Jason Acu�a	http://en.wikipedia.org/wiki/Jason_Acu%F1a
Jason Alexander	http://en.wikipedia.org/wiki/Jason_Alexander
Jason Altmire	http://en.wikipedia.org/wiki/Jason_Altmire
Jason Bateman	http://en.wikipedia.org/wiki/Jason_Bateman
Jason Behr	http://en.wikipedia.org/wiki/Jason_Behr
Jason Biggs	http://en.wikipedia.org/wiki/Jason_Biggs
Jason Chaffetz	http://en.wikipedia.org/wiki/Jason_Chaffetz
Jason Connery	http://en.wikipedia.org/wiki/Jason_Connery
Jason Cook	http://en.wikipedia.org/wiki/Jason_Cook
Jason Donovan	http://en.wikipedia.org/wiki/Jason_Donovan
Jason Evers	http://en.wikipedia.org/wiki/Jason_Evers
Jason Gedrick	http://en.wikipedia.org/wiki/Jason_Gedrick
Jason Giambi	http://en.wikipedia.org/wiki/Jason_Giambi
Jason Gould	http://en.wikipedia.org/wiki/Jason_Gould
Jason Isaacs	http://en.wikipedia.org/wiki/Jason_Isaacs
Jason Jones	http://en.wikipedia.org/wiki/Jason_Jones_(actor)
Jason Kidd	http://en.wikipedia.org/wiki/Jason_Kidd
Jason Lee	http://en.wikipedia.org/wiki/Jason_Lee_(actor)
Jason Lewis	http://en.wikipedia.org/wiki/Jason_Lewis_(actor)
Jason London	http://en.wikipedia.org/wiki/Jason_London
Jason Marsden	http://en.wikipedia.org/wiki/Jason_Marsden
Jason McCartney	http://en.wikipedia.org/wiki/Jason_McCartney_(politician)
Jason Mewes	http://en.wikipedia.org/wiki/Jason_Mewes
Jason Miller	http://en.wikipedia.org/wiki/Jason_Miller_(playwright)
Jason Mraz	http://en.wikipedia.org/wiki/Jason_Mraz
Jason Newsted	http://en.wikipedia.org/wiki/Jason_Newsted
Jason Patric	http://en.wikipedia.org/wiki/Jason_Patric
Jason Priestley	http://en.wikipedia.org/wiki/Jason_Priestley
Jason Ritter	http://en.wikipedia.org/wiki/Jason_Ritter
Jason Robards	http://en.wikipedia.org/wiki/Jason_Robards
Jason Schwartzman	http://en.wikipedia.org/wiki/Jason_Schwartzman
Jason Scott Lee	http://en.wikipedia.org/wiki/Jason_Scott_Lee
Jason Sehorn	http://en.wikipedia.org/wiki/Jason_Sehorn
Jason Statham	http://en.wikipedia.org/wiki/Jason_Statham
Jason Wiles	http://en.wikipedia.org/wiki/Jason_Wiles
Jasper Johns	http://en.wikipedia.org/wiki/Jasper_Johns
Jaume Bartumeu	http://en.wikipedia.org/wiki/Jaume_Bartumeu
Javier Bardem	http://en.wikipedia.org/wiki/Javier_Bardem
Javier P�rez de Cuellar	http://en.wikipedia.org/wiki/Javier_P%E9rez_de_Cuellar
Javier Vel�squez	http://en.wikipedia.org/wiki/Javier_Vel%E1squez
Javy Lopez	http://en.wikipedia.org/wiki/Javy_Lopez
Jawaharlal Nehru	http://en.wikipedia.org/wiki/Jawaharlal_Nehru
Jay Allen	http://en.wikipedia.org/wiki/Jay_Allen
Jay Berwanger	http://en.wikipedia.org/wiki/Jay_Berwanger
Jay Black	http://en.wikipedia.org/wiki/Jay_Black
Jay Cocks	http://en.wikipedia.org/wiki/Jay_Cocks
Jay Garner	http://en.wikipedia.org/wiki/Jay_Garner
Jay Gould	http://en.wikipedia.org/wiki/Jay_Gould
Jay Hernandez	http://en.wikipedia.org/wiki/Jay_Hernandez
Jay Inslee	http://en.wikipedia.org/wiki/Jay_Inslee
Jay Johnston	http://en.wikipedia.org/wiki/Jay_Johnston
Jay Kay	http://en.wikipedia.org/wiki/Jay_Kay
Jay Leno	http://en.wikipedia.org/wiki/Jay_Leno
Jay Macpherson	http://en.wikipedia.org/wiki/Jay_Macpherson
Jay Mohr	http://en.wikipedia.org/wiki/Jay_Mohr
Jay North	http://en.wikipedia.org/wiki/Jay_North
Jay Osmond	http://en.wikipedia.org/wiki/Jay_Osmond
Jay R. Ferguson	http://en.wikipedia.org/wiki/Jay_R._Ferguson
Jay Roach	http://en.wikipedia.org/wiki/Jay_Roach
Jay Rockefeller	http://en.wikipedia.org/wiki/Jay_Rockefeller
Jay Sarno	http://en.wikipedia.org/wiki/Jay_Sarno
Jay Sekulow	http://en.wikipedia.org/wiki/Jay_Sekulow
Jay Silverheels	http://en.wikipedia.org/wiki/Jay_Silverheels
Jay Warren	http://en.wikipedia.org/wiki/Jay_Warren
Jaye Davidson	http://en.wikipedia.org/wiki/Jaye_Davidson
Jayne Brook	http://en.wikipedia.org/wiki/Jayne_Brook
Jayne Kennedy	http://en.wikipedia.org/wiki/Jayne_Kennedy
Jayne Mansfield	http://en.wikipedia.org/wiki/Jayne_Mansfield
Jayne Meadows	http://en.wikipedia.org/wiki/Jayne_Meadows
Jayson Blair	http://en.wikipedia.org/wiki/Jayson_Blair
Jayson Williams	http://en.wikipedia.org/wiki/Jayson_Williams
Jaz Coleman	http://en.wikipedia.org/wiki/Jaz_Coleman
Jean Alesi	http://en.wikipedia.org/wiki/Jean_Alesi
Jean Amila	http://en.wikipedia.org/wiki/Jean_Amila
Jean Anouilh	http://en.wikipedia.org/wiki/Jean_Anouilh
Jean Arp	http://en.wikipedia.org/wiki/Jean_Arp
Jean Arthur	http://en.wikipedia.org/wiki/Jean_Arthur
Jean Baptiste Joseph Fourier	http://en.wikipedia.org/wiki/Jean_Baptiste_Joseph_Fourier
Jean Baudrillard	http://en.wikipedia.org/wiki/Jean_Baudrillard
Jean Bodin	http://en.wikipedia.org/wiki/Jean_Bodin
Jean Buridan	http://en.wikipedia.org/wiki/Jean_Buridan
Jean Charles Tacchella	http://en.wikipedia.org/wiki/Jean-Charles_Tacchella
Jean Chr�tien	http://en.wikipedia.org/wiki/Jean_Chr%E9tien
Jean Cocteau	http://en.wikipedia.org/wiki/Jean_Cocteau
Jean Daurat	http://en.wikipedia.org/wiki/Jean_Daurat
Jean de La Bruy�re	http://en.wikipedia.org/wiki/Jean_de_La_Bruy%E8re
Jean de la Fontaine	http://en.wikipedia.org/wiki/Jean_de_la_Fontaine
Jean Desmarets	http://en.wikipedia.org/wiki/Jean_Desmarets
Jean Eyeghe Ndong	http://en.wikipedia.org/wiki/Jean_Eyeghe_Ndong
Jean Gabin	http://en.wikipedia.org/wiki/Jean_Gabin
Jean Genet	http://en.wikipedia.org/wiki/Jean_Genet
Jean Giraudoux	http://en.wikipedia.org/wiki/Jean_Giraudoux
Jean Hagen	http://en.wikipedia.org/wiki/Jean_Hagen
Jean Hardouin	http://en.wikipedia.org/wiki/Jean_Hardouin
Jean Harlow	http://en.wikipedia.org/wiki/Jean_Harlow
Jean Hersholt	http://en.wikipedia.org/wiki/Jean_Hersholt
Jean I	http://en.wikipedia.org/wiki/John_I_of_France
Jean II	http://en.wikipedia.org/wiki/Jean_II_of_France
Jean Jacques Rousseau	http://en.wikipedia.org/wiki/Jean_Jacques_Rousseau
Jean Jaur�s	http://en.wikipedia.org/wiki/Jean_Jaur%E8s
Jean Kasem	http://en.wikipedia.org/wiki/Jean_Kasem
Jean Langlais	http://en.wikipedia.org/wiki/Jean_Langlais
Jean le Rond d'Alembert	http://en.wikipedia.org/wiki/Jean_le_Rond_d%27Alembert
Jean Louisa Kelly	http://en.wikipedia.org/wiki/Jean_Louisa_Kelly
Jean Marais	http://en.wikipedia.org/wiki/Jean_Marais
Jean Marsh	http://en.wikipedia.org/wiki/Jean_Marsh
Jean Monnet	http://en.wikipedia.org/wiki/Jean_Monnet
Jean Moulin	http://en.wikipedia.org/wiki/Jean_Moulin
Jean Negulesco	http://en.wikipedia.org/wiki/Jean_Negulesco
Jean Nicholas Nicollet	http://en.wikipedia.org/wiki/Jean_Nicholas_Nicollet
Jean Parker	http://en.wikipedia.org/wiki/Jean_Parker
Jean Passerat	http://en.wikipedia.org/wiki/Jean_Passerat
Jean Perrin	http://en.wikipedia.org/wiki/Jean_Perrin
Jean Peters	http://en.wikipedia.org/wiki/Jean_Peters
Jean Piaget	http://en.wikipedia.org/wiki/Jean_Piaget
Jean Racine	http://en.wikipedia.org/wiki/Jean_Racine
Jean Reno	http://en.wikipedia.org/wiki/Jean_Reno
Jean Renoir	http://en.wikipedia.org/wiki/Jean_Renoir
Jean Rhys	http://en.wikipedia.org/wiki/Jean_Rhys
Jean Rochefort	http://en.wikipedia.org/wiki/Jean_Rochefort
Jean Schmidt	http://en.wikipedia.org/wiki/Jean_Schmidt
Jean Seberg	http://en.wikipedia.org/wiki/Jean_Seberg
Jean Senebier	http://en.wikipedia.org/wiki/Jean_Senebier
Jean Shrimpton	http://en.wikipedia.org/wiki/Jean_Shrimpton
Jean Sibelius	http://en.wikipedia.org/wiki/Jean_Sibelius
Jean Simmons	http://en.wikipedia.org/wiki/Jean_Simmons
Jean Smart	http://en.wikipedia.org/wiki/Jean_Smart
Jean Stafford	http://en.wikipedia.org/wiki/Jean_Stafford
Jean Stapleton	http://en.wikipedia.org/wiki/Jean_Stapleton
Jean Toomer	http://en.wikipedia.org/wiki/Jean_Toomer
Jean-Andr� Deluc	http://en.wikipedia.org/wiki/Jean-Andr%E9_Deluc
Jean-Antoine de Ba�f	http://en.wikipedia.org/wiki/Jean-Antoine_de_Ba%EFf
Jean-Antoine Houdon	http://en.wikipedia.org/wiki/Jean-Antoine_Houdon
Jean-Auguste-Dominique Ingres	http://en.wikipedia.org/wiki/Jean-Auguste-Dominique_Ingres
Jean-Baptiste Biot	http://en.wikipedia.org/wiki/Jean-Baptiste_Biot
Jean-Baptiste Colbert	http://en.wikipedia.org/wiki/Jean-Baptiste_Colbert
Jean-Baptiste de Gribeauval	http://en.wikipedia.org/wiki/Jean-Baptiste_de_Gribeauval
Jean-Baptiste Greuze	http://en.wikipedia.org/wiki/Jean-Baptiste_Greuze
Jean-Baptiste Jourdan	http://en.wikipedia.org/wiki/Jean-Baptiste_Jourdan
Jean-Baptiste Lamarck	http://en.wikipedia.org/wiki/Jean-Baptiste_Lamarck
Jean-Baptiste Louvet	http://en.wikipedia.org/wiki/Jean-Baptiste_Louvet
Jean-Baptiste Lully	http://en.wikipedia.org/wiki/Jean-Baptiste_Lully
Jean-Baptiste-Andr� Dumas	http://en.wikipedia.org/wiki/Jean-Baptiste_Dumas
Jean-Baptiste-Joseph Delambre	http://en.wikipedia.org/wiki/Jean-Baptiste-Joseph_Delambre
Jean-Baptiste-Louis Gresset	http://en.wikipedia.org/wiki/Jean-Baptiste-Louis_Gresset
Jean-Benoit Dunckel	http://en.wikipedia.org/wiki/Jean-Benoit_Dunckel
Jean-Bertrand Aristide	http://en.wikipedia.org/wiki/Jean-Bertrand_Aristide
Jean-Charles-Athanase Peltier	http://en.wikipedia.org/wiki/Jean-Charles-Athanase_Peltier
Jean-Claude Duvalier	http://en.wikipedia.org/wiki/Jean-Claude_Duvalier
Jean-Claude Juncker	http://en.wikipedia.org/wiki/Jean-Claude_Juncker
Jean-Claude Killy	http://en.wikipedia.org/wiki/Jean-Claude_Killy
Jean-Claude Pierre-Louis	http://en.wikipedia.org/wiki/Jean-Claude_Pierre-Louis
Jean-Claude Van Damme	http://en.wikipedia.org/wiki/Jean-Claude_Van_Damme
Jeane Dixon	http://en.wikipedia.org/wiki/Jeane_Dixon
Jeane Kirkpatrick	http://en.wikipedia.org/wiki/Jeane_Kirkpatrick
Jean-�tienne Liotard	http://en.wikipedia.org/wiki/Jean-%C9tienne_Liotard
Jeanette MacDonald	http://en.wikipedia.org/wiki/Jeanette_MacDonald
Jeanette Winterson	http://en.wikipedia.org/wiki/Jeanette_Winterson
Jean-Fran�ois Champollion	http://en.wikipedia.org/wiki/Jean-Fran%E7ois_Champollion
Jean-Fran�ois Lyotard	http://en.wikipedia.org/wiki/Jean-Fran%E7ois_Lyotard
Jean-Fran�ois Ntoutoume Emane	http://en.wikipedia.org/wiki/Jean-Fran%E7ois_Ntoutoume_Emane
Jean-Honor� Fragonard	http://en.wikipedia.org/wiki/Jean-Honor%E9_Fragonard
Jeanine Pirro	http://en.wikipedia.org/wiki/Jeanine_Pirro
Jean-Jacques Annaud	http://en.wikipedia.org/wiki/Jean-Jacques_Annaud
Jean-Jacques Rousseau	http://en.wikipedia.org/wiki/Jean-Jacques_Rousseau
Jean-Lambert Tallien	http://en.wikipedia.org/wiki/Jean-Lambert_Tallien
Jean-Leon Gerome	http://en.wikipedia.org/wiki/Jean-Leon_Gerome
Jean-Louis Barrault	http://en.wikipedia.org/wiki/Jean-Louis_Barrault
Jean-Louis Trintignant	http://en.wikipedia.org/wiki/Jean-Louis_Trintignant
Jean-Luc Godard	http://en.wikipedia.org/wiki/Jean-Luc_Godard
Jean-Luc Ponty	http://en.wikipedia.org/wiki/Jean-Luc_Ponty
Jean-Marie Dor�	http://en.wikipedia.org/wiki/Jean-Marie_Dor%E9
Jean-Marie Le Pen	http://en.wikipedia.org/wiki/Jean-Marie_Le_Pen
Jean-Marie Lehn	http://en.wikipedia.org/wiki/Jean-Marie_Lehn
Jean-Marie Messier	http://en.wikipedia.org/wiki/Jean-Marie_Messier
Jean-Marie Roland	http://en.wikipedia.org/wiki/Jean-Marie_Roland
Jean-Max Bellerive	http://en.wikipedia.org/wiki/Jean-Max_Bellerive
Jean-Michel Basquiat	http://en.wikipedia.org/wiki/Jean-Michel_Basquiat
Jean-Michel Jarre	http://en.wikipedia.org/wiki/Jean-Michel_Jarre
Jeanne Calment	http://en.wikipedia.org/wiki/Jeanne_Calment
Jeanne Crain	http://en.wikipedia.org/wiki/Jeanne_Crain
Jeanne Moreau	http://en.wikipedia.org/wiki/Jeanne_Moreau
Jeanne Shaheen	http://en.wikipedia.org/wiki/Jeanne_Shaheen
Jeanne Tripplehorn	http://en.wikipedia.org/wiki/Jeanne_Tripplehorn
Jeanne-Marie Roland	http://en.wikipedia.org/wiki/Jeanne-Marie_Roland
Jean-Paul Belmondo	http://en.wikipedia.org/wiki/Jean-Paul_Belmondo
Jean-Paul Gaultier	http://en.wikipedia.org/wiki/Jean-Paul_Gaultier
Jean-Paul Marat	http://en.wikipedia.org/wiki/Jean-Paul_Marat
Jean-Paul Proust	http://en.wikipedia.org/wiki/Jean-Paul_Proust
Jean-Paul Sartre	http://en.wikipedia.org/wiki/Jean-Paul_Sartre
Jean-Philippe Rameau	http://en.wikipedia.org/wiki/Jean-Philippe_Rameau
Jean-Pierre Boyer	http://en.wikipedia.org/wiki/Jean-Pierre_Boyer
Jean-Pierre Cassel	http://en.wikipedia.org/wiki/Jean-Pierre_Cassel
Jean-Pierre Jeunet	http://en.wikipedia.org/wiki/Jean-Pierre_Jeunet
Jean-Pierre Mocky	http://en.wikipedia.org/wiki/Jean-Pierre_Mocky
Jean-Pierre Raffarin	http://en.wikipedia.org/wiki/Jean-Pierre_Raffarin
Jean-Sylvain Bailly	http://en.wikipedia.org/wiki/Jean-Sylvain_Bailly
Jeb Bradley	http://en.wikipedia.org/wiki/Jeb_Bradley
Jeb Bush	http://en.wikipedia.org/wiki/Jeb_Bush
Jeb Bush	http://en.wikipedia.org/wiki/Jeb_Bush
Jeb Hensarling	http://en.wikipedia.org/wiki/Jeb_Hensarling
Jeb Magruder	http://en.wikipedia.org/wiki/Jeb_Magruder
Jeb Stuart	http://en.wikipedia.org/wiki/Jeb_Stuart
Jebby Bush	http://en.wikipedia.org/wiki/Jebby_Bush
Jef Raskin	http://en.wikipedia.org/wiki/Jef_Raskin
Jeff Altman	http://en.wikipedia.org/wiki/Jeff_Altman
Jeff Ament	http://en.wikipedia.org/wiki/Jeff_Ament
Jeff Beck	http://en.wikipedia.org/wiki/Jeff_Beck
Jeff Bezos	http://en.wikipedia.org/wiki/Jeff_Bezos
Jeff Bingaman	http://en.wikipedia.org/wiki/Jeff_Bingaman
Jeff Bingaman	http://en.wikipedia.org/wiki/Jeff_Bingaman
Jeff Bridges	http://en.wikipedia.org/wiki/Jeff_Bridges
Jeff Buckley	http://en.wikipedia.org/wiki/Jeff_Buckley
Jeff Chandler	http://en.wikipedia.org/wiki/Jeff_Chandler_(actor)
Jeff Cohen	http://en.wikipedia.org/wiki/Jeff_Cohen_(media_critic)
Jeff Conaway	http://en.wikipedia.org/wiki/Jeff_Conaway
Jeff Daniels	http://en.wikipedia.org/wiki/Jeff_Daniels
Jeff Dowd	http://en.wikipedia.org/wiki/Jeff_Dowd
Jeff Fahey	http://en.wikipedia.org/wiki/Jeff_Fahey
Jeff Flake	http://en.wikipedia.org/wiki/Jeff_Flake
Jeff Fortenberry	http://en.wikipedia.org/wiki/Jeff_Fortenberry
Jeff Foxworthy	http://en.wikipedia.org/wiki/Jeff_Foxworthy
Jeff Gannon	http://en.wikipedia.org/wiki/Jeff_Gannon
Jeff Garcia	http://en.wikipedia.org/wiki/Jeff_Garcia
Jeff Goldblum	http://en.wikipedia.org/wiki/Jeff_Goldblum
Jeff Gordon	http://en.wikipedia.org/wiki/Jeff_Gordon
Jeff Greenfield	http://en.wikipedia.org/wiki/Jeff_Greenfield
Jeff Habay	http://en.wikipedia.org/wiki/Jeff_Habay
Jeff Hanneman	http://en.wikipedia.org/wiki/Jeff_Hanneman
Jeff Hoffman	http://en.wikipedia.org/wiki/Jeff_Hoffman
Jeff Koons	http://en.wikipedia.org/wiki/Jeff_Koons
Jeff Lieberman	http://en.wikipedia.org/wiki/Jeff_Lieberman
Jeff Lynne	http://en.wikipedia.org/wiki/Jeff_Lynne
Jeff MacNelly	http://en.wikipedia.org/wiki/Jeff_MacNelly
Jeff Merkley	http://en.wikipedia.org/wiki/Jeff_Merkley
Jeff Miller	http://en.wikipedia.org/wiki/Jeff_Miller
Jeff Probst	http://en.wikipedia.org/wiki/Jeff_Probst
Jeff Sessions	http://en.wikipedia.org/wiki/Jeff_Sessions
Jeff Skoll	http://en.wikipedia.org/wiki/Jeff_Skoll
Jeff Smith	http://en.wikipedia.org/wiki/Jeff_Smith_(TV_personality)
Jeff Tremaine	http://en.wikipedia.org/wiki/Jeff_Tremaine
Jeff Tweedy	http://en.wikipedia.org/wiki/Jeff_Tweedy
Jeff Vandermeer	http://en.wikipedia.org/wiki/Jeff_Vandermeer
Jefferson Davis	http://en.wikipedia.org/wiki/Jefferson_Davis
Jefferson Hack	http://en.wikipedia.org/wiki/Jefferson_Hack
Jeffrey A. Joerres	http://en.wikipedia.org/wiki/Jeffrey_A._Joerres
Jeffrey Cohelan	http://en.wikipedia.org/wiki/Jeffrey_Cohelan
Jeffrey Combs	http://en.wikipedia.org/wiki/Jeffrey_Combs
Jeffrey Dahmer	http://en.wikipedia.org/wiki/Jeffrey_Dahmer
Jeffrey Eugenides	http://en.wikipedia.org/wiki/Jeffrey_Eugenides
Jeffrey Hunter	http://en.wikipedia.org/wiki/Jeffrey_Hunter
Jeffrey Jones	http://en.wikipedia.org/wiki/Jeffrey_Jones
Jeffrey Katzenberg	http://en.wikipedia.org/wiki/Jeffrey_Katzenberg
Jeffrey Loria	http://en.wikipedia.org/wiki/Jeffrey_Loria
Jeffrey M. Donaldson	http://en.wikipedia.org/wiki/Jeffrey_Donaldson
Jeffrey Osborne	http://en.wikipedia.org/wiki/Jeffrey_Osborne
Jeffrey R. Immelt	http://en.wikipedia.org/wiki/Jeffrey_R._Immelt
Jeffrey Sachs	http://en.wikipedia.org/wiki/Jeffrey_Sachs
Jeffrey Skilling	http://en.wikipedia.org/wiki/Jeffrey_Skilling
Jeffrey Tambor	http://en.wikipedia.org/wiki/Jeffrey_Tambor
Jeffrey Wright	http://en.wikipedia.org/wiki/Jeffrey_Wright_(actor)
Jello Biafra	http://en.wikipedia.org/wiki/Jello_Biafra
Jelly Roll Morton	http://en.wikipedia.org/wiki/Jelly_Roll_Morton
Jena Malone	http://en.wikipedia.org/wiki/Jena_Malone
Jenette Goldstein	http://en.wikipedia.org/wiki/Jenette_Goldstein
Jenifer Lewis	http://en.wikipedia.org/wiki/Jenifer_Lewis
Jenilee Harrison	http://en.wikipedia.org/wiki/Jenilee_Harrison
Jenna Bush	http://en.wikipedia.org/wiki/Jenna_Bush
Jenna Elfman	http://en.wikipedia.org/wiki/Jenna_Elfman
Jenna Jameson	http://en.wikipedia.org/wiki/Jenna_Jameson
Jenna von Oy	http://en.wikipedia.org/wiki/Jenna_von_Oy
Jennette Bradley	http://en.wikipedia.org/wiki/Jennette_Bradley
Jennie Garth	http://en.wikipedia.org/wiki/Jennie_Garth
Jennifer 8. Lee	http://en.wikipedia.org/wiki/Jennifer_8._Lee
Jennifer Aniston	http://en.wikipedia.org/wiki/Jennifer_Aniston
Jennifer Beals	http://en.wikipedia.org/wiki/Jennifer_Beals
Jennifer Capriati	http://en.wikipedia.org/wiki/Jennifer_Capriati
Jennifer Connelly	http://en.wikipedia.org/wiki/Jennifer_Connelly
Jennifer Coolidge	http://en.wikipedia.org/wiki/Jennifer_Coolidge
Jennifer Dunn	http://en.wikipedia.org/wiki/Jennifer_Dunn
Jennifer Ehle	http://en.wikipedia.org/wiki/Jennifer_Ehle
Jennifer Esposito	http://en.wikipedia.org/wiki/Jennifer_Esposito
Jennifer Finch	http://en.wikipedia.org/wiki/Jennifer_Finch
Jennifer Freeman	http://en.wikipedia.org/wiki/Jennifer_Freeman
Jennifer Garner	http://en.wikipedia.org/wiki/Jennifer_Garner
Jennifer Granholm	http://en.wikipedia.org/wiki/Jennifer_Granholm
Jennifer Granholm	http://en.wikipedia.org/wiki/Jennifer_Granholm
Jennifer Granick	http://en.wikipedia.org/wiki/Jennifer_Granick
Jennifer Grey	http://en.wikipedia.org/wiki/Jennifer_Grey
Jennifer Jason Leigh	http://en.wikipedia.org/wiki/Jennifer_Jason_Leigh
Jennifer Jones	http://en.wikipedia.org/wiki/Jennifer_Jones
Jennifer Lopez	http://en.wikipedia.org/wiki/Jennifer_Lopez
Jennifer Love Hewitt	http://en.wikipedia.org/wiki/Jennifer_Love_Hewitt
Jennifer O'Neill	http://en.wikipedia.org/wiki/Jennifer_O%27Neill
Jennifer Saunders	http://en.wikipedia.org/wiki/Jennifer_Saunders
Jennifer Tilly	http://en.wikipedia.org/wiki/Jennifer_Tilly
Jennifer Vanderbes	http://en.wikipedia.org/wiki/Jennifer_Vanderbes
Jenny Agutter	http://en.wikipedia.org/wiki/Jenny_Agutter
Jenny Chapman	http://en.wikipedia.org/wiki/Jenny_Chapman
Jenny Jones	http://en.wikipedia.org/wiki/Jenny_Jones_(presenter)
Jenny Lewis	http://en.wikipedia.org/wiki/Jenny_Lewis
Jenny McCarthy	http://en.wikipedia.org/wiki/Jenny_McCarthy
Jenny Shimizu	http://en.wikipedia.org/wiki/Jenny_Shimizu
Jenny Willott	http://en.wikipedia.org/wiki/Jenny_Willott
Jens Albinus	http://en.wikipedia.org/wiki/Jens_Albinus
Jens B�hrnsen	http://en.wikipedia.org/wiki/Jens_B%F6hrnsen
Jens C. Skou	http://en.wikipedia.org/wiki/Jens_C._Skou
Jens Peter Jacobsen	http://en.wikipedia.org/wiki/Jens_Peter_Jacobsen
Jens Stoltenberg	http://en.wikipedia.org/wiki/Jens_Stoltenberg
Jensen Ackles	http://en.wikipedia.org/wiki/Jensen_Ackles
Jerald F. ter Horst	http://en.wikipedia.org/wiki/Jerald_terHorst
Jeremiah A. Denton Jr.	http://en.wikipedia.org/wiki/Jeremiah_Denton
Jeremiah Horrocks	http://en.wikipedia.org/wiki/Jeremiah_Horrocks
Jeremy Akerman	http://en.wikipedia.org/wiki/Jeremy_Akerman
Jeremy Bentham	http://en.wikipedia.org/wiki/Jeremy_Bentham
Jeremy Brett	http://en.wikipedia.org/wiki/Jeremy_Brett
Jeremy Browne	http://en.wikipedia.org/wiki/Jeremy_Browne
Jeremy Bulloch	http://en.wikipedia.org/wiki/Jeremy_Bulloch
Jeremy Corbyn	http://en.wikipedia.org/wiki/Jeremy_Corbyn
Jeremy Hunt	http://en.wikipedia.org/wiki/Jeremy_Hunt_(politician)
Jeremy Irons	http://en.wikipedia.org/wiki/Jeremy_Irons
Jeremy Jackson	http://en.wikipedia.org/wiki/Jeremy_Jackson
Jeremy Lefroy	http://en.wikipedia.org/wiki/Jeremy_Lefroy
Jeremy Leven	http://en.wikipedia.org/wiki/Jeremy_Leven
Jeremy London	http://en.wikipedia.org/wiki/Jeremy_London
Jeremy Miller	http://en.wikipedia.org/wiki/Jeremy_Miller
Jeremy Northam	http://en.wikipedia.org/wiki/Jeremy_Northam
Jeremy Piven	http://en.wikipedia.org/wiki/Jeremy_Piven
Jeremy Rifkin	http://en.wikipedia.org/wiki/Jeremy_Rifkin
Jeremy Sisto	http://en.wikipedia.org/wiki/Jeremy_Sisto
Jeremy Sumpter	http://en.wikipedia.org/wiki/Jeremy_Sumpter
Jeremy Taylor	http://en.wikipedia.org/wiki/Jeremy_Taylor
Jeremy Wright	http://en.wikipedia.org/wiki/Jeremy_Wright_(politician)
Jeri Ryan	http://en.wikipedia.org/wiki/Jeri_Ryan
Jermaine Dupri	http://en.wikipedia.org/wiki/Jermaine_Dupri
Jermaine Jackson	http://en.wikipedia.org/wiki/Jermaine_Jackson
Jerome Alden	http://en.wikipedia.org/wiki/Jerome_Alden
Jerome Bettis	http://en.wikipedia.org/wiki/Jerome_Bettis
Jerome Corsi	http://en.wikipedia.org/wiki/Jerome_Corsi
Jerome I. Friedman	http://en.wikipedia.org/wiki/Jerome_I._Friedman
Jerome K. Jerome	http://en.wikipedia.org/wiki/Jerome_K._Jerome
Jerome Karle	http://en.wikipedia.org/wiki/Jerome_Karle
Jerome Lawrence	http://en.wikipedia.org/wiki/Jerome_Lawrence
Jerome Robbins	http://en.wikipedia.org/wiki/Jerome_Robbins
Jerrold Nadler	http://en.wikipedia.org/wiki/Jerrold_Nadler
Jerry A. Grundhofer	http://en.wikipedia.org/wiki/Jerry_Grundhofer
Jerry Bailey	http://en.wikipedia.org/wiki/Jerry_Bailey
Jerry Boykin	http://en.wikipedia.org/wiki/William_G._Boykin
Jerry Brown	http://en.wikipedia.org/wiki/Jerry_Brown
Jerry Bruckheimer	http://en.wikipedia.org/wiki/Jerry_Bruckheimer
Jerry Butler	http://en.wikipedia.org/wiki/Jerry_Butler_(singer)
Jerry Cantrell	http://en.wikipedia.org/wiki/Jerry_Cantrell
Jerry Costello	http://en.wikipedia.org/wiki/Jerry_Costello
Jerry Doyle	http://en.wikipedia.org/wiki/Jerry_Doyle_(radio_host)
Jerry Falwell	http://en.wikipedia.org/wiki/Jerry_Falwell
Jerry Garcia	http://en.wikipedia.org/wiki/Jerry_Garcia
Jerry Goldsmith	http://en.wikipedia.org/wiki/Jerry_Goldsmith
Jerry Greenfield	http://en.wikipedia.org/wiki/Jerry_Greenfield
Jerry Hall	http://en.wikipedia.org/wiki/Jerry_Hall
Jerry Harrison	http://en.wikipedia.org/wiki/Jerry_Harrison
Jerry Jeff Walker	http://en.wikipedia.org/wiki/Jerry_Jeff_Walker
Jerry Jones	http://en.wikipedia.org/wiki/Jerry_Jones
Jerry Juhl	http://en.wikipedia.org/wiki/Jerry_Juhl
Jerry Kleczka	http://en.wikipedia.org/wiki/Jerry_Kleczka
Jerry Lawler	http://en.wikipedia.org/wiki/Jerry_Lawler
Jerry Lee Lewis	http://en.wikipedia.org/wiki/Jerry_Lee_Lewis
Jerry Leiber	http://en.wikipedia.org/wiki/Jerry_Leiber
Jerry Levin	http://en.wikipedia.org/wiki/Jerry_Levin
Jerry Lewis	http://en.wikipedia.org/wiki/Jerry_Lewis
Jerry Lewis	http://en.wikipedia.org/wiki/Jerry_Lewis_(politician)
Jerry Lewis	http://en.wikipedia.org/wiki/Jerry_Lewis_(politician)
Jerry Marotta	http://en.wikipedia.org/wiki/Jerry_Marotta
Jerry Mathers	http://en.wikipedia.org/wiki/Jerry_Mathers
Jerry McNerney	http://en.wikipedia.org/wiki/Jerry_McNerney
Jerry Moran	http://en.wikipedia.org/wiki/Jerry_Moran
Jerry Moss	http://en.wikipedia.org/wiki/Jerry_Moss
Jerry Nachman	http://en.wikipedia.org/wiki/Jerry_Nachman
Jerry O'Connell	http://en.wikipedia.org/wiki/Jerry_O%27Connell
Jerry Only	http://en.wikipedia.org/wiki/Jerry_Only
Jerry Orbach	http://en.wikipedia.org/wiki/Jerry_Orbach
Jerry Perenchio	http://en.wikipedia.org/wiki/Jerry_Perenchio
Jerry Pournelle	http://en.wikipedia.org/wiki/Jerry_Pournelle
Jerry Reed	http://en.wikipedia.org/wiki/Jerry_Reed
Jerry Rice	http://en.wikipedia.org/wiki/Jerry_Rice
Jerry Rubin	http://en.wikipedia.org/wiki/Jerry_Rubin
Jerry Seinfeld	http://en.wikipedia.org/wiki/Jerry_Seinfeld
Jerry Springer	http://en.wikipedia.org/wiki/Jerry_Springer
Jerry Stahl	http://en.wikipedia.org/wiki/Jerry_Stahl
Jerry Stiller	http://en.wikipedia.org/wiki/Jerry_Stiller
Jerry Tarkanian	http://en.wikipedia.org/wiki/Jerry_Tarkanian
Jerry Vale	http://en.wikipedia.org/wiki/Jerry_Vale
Jerry Van Dyke	http://en.wikipedia.org/wiki/Jerry_Van_Dyke
Jerry Weller	http://en.wikipedia.org/wiki/Jerry_Weller
Jerry Yang	http://en.wikipedia.org/wiki/Jerry_Yang_(entrepreneur)
Jerry Zucker	http://en.wikipedia.org/wiki/Jerry_Zucker_(film_director)
Jeru the Damaja	http://en.wikipedia.org/wiki/Jeru_the_Damaja
Jerzy Kosinski	http://en.wikipedia.org/wiki/Jerzy_Kosinski
Jerzy Popieluszko	http://en.wikipedia.org/wiki/Jerzy_Popieluszko
Jessamyn West	http://en.wikipedia.org/wiki/Jessamyn_West_(writer)
Jesse Bradford	http://en.wikipedia.org/wiki/Jesse_Bradford
Jesse Brown	http://en.wikipedia.org/wiki/Jesse_Brown
Jesse H. Jones	http://en.wikipedia.org/wiki/Jesse_H._Jones
Jesse Helms	http://en.wikipedia.org/wiki/Jesse_Helms
Jesse Helms	http://en.wikipedia.org/wiki/Jesse_Helms
Jesse Jackson	http://en.wikipedia.org/wiki/Jesse_Jackson
Jesse Jackson, Jr.	http://en.wikipedia.org/wiki/Jesse_Jackson%2C_Jr.
Jesse James	http://en.wikipedia.org/wiki/Jesse_James_(customizer)
Jesse James	http://en.wikipedia.org/wiki/Jesse_James
Jesse L. Martin	http://en.wikipedia.org/wiki/Jesse_L._Martin
Jesse Martin Combs	http://en.wikipedia.org/wiki/Jesse_Martin_Combs
Jesse McCartney	http://en.wikipedia.org/wiki/Jesse_McCartney
Jesse Metcalfe	http://en.wikipedia.org/wiki/Jesse_Metcalfe
Jesse Norman	http://en.wikipedia.org/wiki/Jesse_Norman
Jesse Owens	http://en.wikipedia.org/wiki/Jesse_Owens
Jesse Spencer	http://en.wikipedia.org/wiki/Jesse_Spencer
Jesse Unruh	http://en.wikipedia.org/wiki/Jesse_Unruh
Jesse Ventura	http://en.wikipedia.org/wiki/Jesse_Ventura
Jessi Colter	http://en.wikipedia.org/wiki/Jessi_Colter
Jessica Alba	http://en.wikipedia.org/wiki/Jessica_Alba
Jessica Biel	http://en.wikipedia.org/wiki/Jessica_Biel
Jessica Cutler	http://en.wikipedia.org/wiki/Jessica_Cutler
Jessica Hagedorn	http://en.wikipedia.org/wiki/Jessica_Hagedorn
Jessica Hahn	http://en.wikipedia.org/wiki/Jessica_Hahn
Jessica Harper	http://en.wikipedia.org/wiki/Jessica_Harper
Jessica Lange	http://en.wikipedia.org/wiki/Jessica_Lange
Jessica Lee	http://en.wikipedia.org/wiki/Jessica_Lee_(politician)
Jessica Lynch	http://en.wikipedia.org/wiki/Jessica_Lynch
Jessica Mitford	http://en.wikipedia.org/wiki/Jessica_Mitford
Jessica Morden	http://en.wikipedia.org/wiki/Jessica_Morden
Jessica Savitch	http://en.wikipedia.org/wiki/Jessica_Savitch
Jessica Simpson	http://en.wikipedia.org/wiki/Jessica_Simpson
Jessica Tandy	http://en.wikipedia.org/wiki/Jessica_Tandy
Jessica Walter	http://en.wikipedia.org/wiki/Jessica_Walter
Jessie Matthews	http://en.wikipedia.org/wiki/Jessie_Matthews
Jessie Redmon Fauset	http://en.wikipedia.org/wiki/Jessie_Redmon_Fauset
Jessie Wilcox Smith	http://en.wikipedia.org/wiki/Jessie_Wilcox_Smith
Jessye Norman	http://en.wikipedia.org/wiki/Jessye_Norman
Jesus Christ	http://en.wikipedia.org/wiki/Jesus_Christ
Jet Li	http://en.wikipedia.org/wiki/Jet_Li
Jethro Tull	http://en.wikipedia.org/wiki/Jethro_Tull_(agriculturist)
Jhonen Vasquez	http://en.wikipedia.org/wiki/Jhonen_Vasquez
Jhumpa Lahiri	http://en.wikipedia.org/wiki/Jhumpa_Lahiri
Jiang Zemin	http://en.wikipedia.org/wiki/Jiang_Zemin
Jigme Singye Wangchuck	http://en.wikipedia.org/wiki/Jigme_Singye_Wangchuck
Jigme Thinley	http://en.wikipedia.org/wiki/Jigme_Thinley
Jill Bennett	http://en.wikipedia.org/wiki/Jill_Bennett_(British_actress)
Jill Clayburgh	http://en.wikipedia.org/wiki/Jill_Clayburgh
Jill Goodacre	http://en.wikipedia.org/wiki/Jill_Goodacre
Jill Hennessy	http://en.wikipedia.org/wiki/Jill_Hennessy
Jill Ireland	http://en.wikipedia.org/wiki/Jill_Ireland
Jill Scott	http://en.wikipedia.org/wiki/Jill_Scott
Jill St. John	http://en.wikipedia.org/wiki/Jill_St._John
Jill Talley	http://en.wikipedia.org/wiki/Jill_Talley
Jillian Parry	http://en.wikipedia.org/wiki/Jillian_Parry
Jim Backus	http://en.wikipedia.org/wiki/Jim_Backus
Jim Bakker	http://en.wikipedia.org/wiki/Jim_Bakker
Jim Barksdale	http://en.wikipedia.org/wiki/Jim_Barksdale
Jim Bates	http://en.wikipedia.org/wiki/Jim_Bates
Jim Beaver	http://en.wikipedia.org/wiki/Jim_Beaver
Jim Bell	http://en.wikipedia.org/wiki/Jim_Bell
Jim Belushi	http://en.wikipedia.org/wiki/Jim_Belushi
Jim Broadbent	http://en.wikipedia.org/wiki/Jim_Broadbent
Jim Brown	http://en.wikipedia.org/wiki/Jim_Brown
Jim Bunning	http://en.wikipedia.org/wiki/Jim_Bunning
Jim Byrnes	http://en.wikipedia.org/wiki/Jim_Byrnes_(actor)
Jim Cantalupo	http://en.wikipedia.org/wiki/Jim_Cantalupo
Jim Carrey	http://en.wikipedia.org/wiki/Jim_Carrey
Jim Chapman	http://en.wikipedia.org/wiki/Jim_Chapman
Jim Clyburn	http://en.wikipedia.org/wiki/Jim_Clyburn
Jim Cooper	http://en.wikipedia.org/wiki/Jim_Cooper
Jim Cooper	http://en.wikipedia.org/wiki/Jim_Cooper
Jim Costa	http://en.wikipedia.org/wiki/Jim_Costa
Jim Courier	http://en.wikipedia.org/wiki/Jim_Courier
Jim Courter	http://en.wikipedia.org/wiki/Jim_Courter
Jim Cramer	http://en.wikipedia.org/wiki/Jim_Cramer
Jim Croce	http://en.wikipedia.org/wiki/Jim_Croce
Jim Cunningham	http://en.wikipedia.org/wiki/Jim_Cunningham_(UK_politician)
Jim Dale	http://en.wikipedia.org/wiki/Jim_Dale
Jim Davis	http://en.wikipedia.org/wiki/Jim_Davis_(cartoonist)
Jim Davis	http://en.wikipedia.org/wiki/Jim_Davis_(politician)
Jim Davis	http://en.wikipedia.org/wiki/Jim_Davis_(actor)
Jim DeMint	http://en.wikipedia.org/wiki/Jim_DeMint
Jim Dobbin	http://en.wikipedia.org/wiki/Jim_Dobbin
Jim Douglas	http://en.wikipedia.org/wiki/Jim_Douglas
Jim Dowd	http://en.wikipedia.org/wiki/Jim_Dowd_(politician)
Jim Doyle	http://en.wikipedia.org/wiki/Jim_Doyle
Jim Ellis	http://en.wikipedia.org/wiki/Jim_Ellis_(computing)
Jim Exon	http://en.wikipedia.org/wiki/Jim_Exon
Jim Fisk	http://en.wikipedia.org/wiki/James_Fisk_(financier)
Jim Fitzpatrick	http://en.wikipedia.org/wiki/Jim_Fitzpatrick_(politician)
Jim Fowler	http://en.wikipedia.org/wiki/Jim_Fowler
Jim Garrison	http://en.wikipedia.org/wiki/Jim_Garrison
Jim Gerlach	http://en.wikipedia.org/wiki/Jim_Gerlach
Jim Gibbons	http://en.wikipedia.org/wiki/Jim_Gibbons_(U.S._politician)
Jim Gilmore	http://en.wikipedia.org/wiki/Jim_Gilmore
Jim Goad	http://en.wikipedia.org/wiki/Jim_Goad
Jim Guy Tucker	http://en.wikipedia.org/wiki/Jim_Guy_Tucker
Jim Henson	http://en.wikipedia.org/wiki/Jim_Henson
Jim Hightower	http://en.wikipedia.org/wiki/Jim_Hightower
Jim Himes	http://en.wikipedia.org/wiki/Jim_Himes
Jim Hoagland	http://en.wikipedia.org/wiki/Jim_Hoagland
Jim Hodges	http://en.wikipedia.org/wiki/Jim_Hodges
Jim Hood	http://en.wikipedia.org/wiki/Jim_Hood
Jim Hutton	http://en.wikipedia.org/wiki/Jim_Hutton
Jim J. Bullock	http://en.wikipedia.org/wiki/Jim_J._Bullock
Jim Jarmusch	http://en.wikipedia.org/wiki/Jim_Jarmusch
Jim Jeffords	http://en.wikipedia.org/wiki/Jim_Jeffords
Jim Jones	http://en.wikipedia.org/wiki/Jim_Jones
Jim Jordan	http://en.wikipedia.org/wiki/Jim_Jordan_(Ohio_politician)
Jim Kaat	http://en.wikipedia.org/wiki/Jim_Kaat
Jim Kelly	http://en.wikipedia.org/wiki/Jim_Kelly
Jim Kerr	http://en.wikipedia.org/wiki/Jim_Kerr
Jim Kolbe	http://en.wikipedia.org/wiki/Jim_Kolbe
Jim Kolbe	http://en.wikipedia.org/wiki/Jim_Kolbe
Jim Lange	http://en.wikipedia.org/wiki/Jim_Lange
Jim Langevin	http://en.wikipedia.org/wiki/Jim_Langevin
Jim Leach	http://en.wikipedia.org/wiki/Jim_Leach
Jim Lehrer	http://en.wikipedia.org/wiki/Jim_Lehrer
Jim Lovell	http://en.wikipedia.org/wiki/Jim_Lovell
Jim Marshall	http://en.wikipedia.org/wiki/Jim_Marshall_(Georgia_politician)
Jim Marurai	http://en.wikipedia.org/wiki/Jim_Marurai
Jim Matheson	http://en.wikipedia.org/wiki/Jim_Matheson
Jim McCrery	http://en.wikipedia.org/wiki/Jim_McCrery
Jim McGovern	http://en.wikipedia.org/wiki/Jim_McGovern
Jim McKay	http://en.wikipedia.org/wiki/Jim_McKay
Jim McMahon	http://en.wikipedia.org/wiki/Jim_McMahon
Jim Messina	http://en.wikipedia.org/wiki/Jim_Messina_(musician)
Jim Mitchell	http://en.wikipedia.org/wiki/Mitchell_brothers
Jim Moody	http://en.wikipedia.org/wiki/Jim_Moody
Jim Moran	http://en.wikipedia.org/wiki/Jim_Moran
Jim Morrison	http://en.wikipedia.org/wiki/Jim_Morrison
Jim Murphy	http://en.wikipedia.org/wiki/Jim_Murphy
Jim Nabors	http://en.wikipedia.org/wiki/Jim_Nabors
Jim Nicholson	http://en.wikipedia.org/wiki/Jim_Nicholson_(U.S._politician)
Jim Norton	http://en.wikipedia.org/wiki/Jim_Norton_(comedian)
Jim Nussle	http://en.wikipedia.org/wiki/Jim_Nussle
Jim Olin	http://en.wikipedia.org/wiki/Jim_Olin
Jim O'Rourke	http://en.wikipedia.org/wiki/Jim_O'Rourke_(musician)
Jim Otto	http://en.wikipedia.org/wiki/Jim_Otto
Jim Palmer	http://en.wikipedia.org/wiki/Jim_Palmer
Jim Pinkerton	http://en.wikipedia.org/wiki/Jim_Pinkerton
Jim Plunkett	http://en.wikipedia.org/wiki/Jim_Plunkett
Jim Ramstad	http://en.wikipedia.org/wiki/Jim_Ramstad
Jim Reeves	http://en.wikipedia.org/wiki/Jim_Reeves
Jim Risch	http://en.wikipedia.org/wiki/Jim_Risch
Jim Rogan	http://en.wikipedia.org/wiki/Jim_Rogan
Jim Rome	http://en.wikipedia.org/wiki/Jim_Rome
Jim Romenesko	http://en.wikipedia.org/wiki/Jim_Romenesko
Jim Rose	http://en.wikipedia.org/wiki/Jim_Rose
Jim Ross Lightfoot	http://en.wikipedia.org/wiki/Jim_Ross_Lightfoot
Jim Ryun	http://en.wikipedia.org/wiki/Jim_Ryun
Jim Sasser	http://en.wikipedia.org/wiki/Jim_Sasser
Jim Sasser	http://en.wikipedia.org/wiki/Jim_Sasser
Jim Saxton	http://en.wikipedia.org/wiki/Jim_Saxton
Jim Sensenbrenner	http://en.wikipedia.org/wiki/Jim_Sensenbrenner
Jim Shannon	http://en.wikipedia.org/wiki/Jim_Shannon
Jim Sheridan	http://en.wikipedia.org/wiki/Jim_Sheridan_(politician)
Jim Skinner	http://en.wikipedia.org/wiki/Jim_Skinner
Jim Slattery	http://en.wikipedia.org/wiki/Jim_Slattery
Jim South	http://en.wikipedia.org/wiki/Jim_South
Jim Talent	http://en.wikipedia.org/wiki/Jim_Talent
Jim Thome	http://en.wikipedia.org/wiki/Jim_Thome
Jim Thompson	http://en.wikipedia.org/wiki/Jim_Thompson_(writer)
Jim Thorpe	http://en.wikipedia.org/wiki/Jim_Thorpe
Jim Turner	http://en.wikipedia.org/wiki/Jim_Turner_(comedian)
Jim Turner	http://en.wikipedia.org/wiki/Jim_Turner_(politician)
Jim Varney	http://en.wikipedia.org/wiki/Jim_Varney
Jim Walsh	http://en.wikipedia.org/wiki/James_T._Walsh
Jim Walton	http://en.wikipedia.org/wiki/Jim_Walton
Jim Webb	http://en.wikipedia.org/wiki/Jim_Webb
Jim Woodring	http://en.wikipedia.org/wiki/Jim_Woodring
Jim Wright	http://en.wikipedia.org/wiki/Jim_Wright
Jim Wright	http://en.wikipedia.org/wiki/Jim_Wright
Jimbo Wales	http://en.wikipedia.org/wiki/Jimbo_Wales
Jimi Hendrix	http://en.wikipedia.org/wiki/Jimi_Hendrix
Jimmie Davis	http://en.wikipedia.org/wiki/Jimmie_Davis
Jimmie Foxx	http://en.wikipedia.org/wiki/Jimmie_Foxx
Jimmie Walker	http://en.wikipedia.org/wiki/Jimmie_Walker
Jimmy Breslin	http://en.wikipedia.org/wiki/Jimmy_Breslin
Jimmy Buffett	http://en.wikipedia.org/wiki/Jimmy_Buffett
Jimmy Carl Black	http://en.wikipedia.org/wiki/Jimmy_Carl_Black
Jimmy Carter	http://en.wikipedia.org/wiki/Jimmy_Carter
Jimmy Castor	http://en.wikipedia.org/wiki/Jimmy_Castor
Jimmy Chamberlin	http://en.wikipedia.org/wiki/Jimmy_Chamberlin
Jimmy Cliff	http://en.wikipedia.org/wiki/Jimmy_Cliff
Jimmy Connors	http://en.wikipedia.org/wiki/Jimmy_Connors
Jimmy Dodd	http://en.wikipedia.org/wiki/Jimmy_Dodd
Jimmy Dorsey	http://en.wikipedia.org/wiki/Jimmy_Dorsey
Jimmy Durante	http://en.wikipedia.org/wiki/Jimmy_Durante
Jimmy Fallon	http://en.wikipedia.org/wiki/Jimmy_Fallon
Jimmy Greaves	http://en.wikipedia.org/wiki/Jimmy_Greaves
Jimmy Hanley	http://en.wikipedia.org/wiki/Jimmy_Hanley
Jimmy Hoffa	http://en.wikipedia.org/wiki/Jimmy_Hoffa
Jimmy Johnstone	http://en.wikipedia.org/wiki/Jimmy_Johnstone
Jimmy Kimmel	http://en.wikipedia.org/wiki/Jimmy_Kimmel
Jimmy McNichol	http://en.wikipedia.org/wiki/Jimmy_McNichol
Jimmy Osmond	http://en.wikipedia.org/wiki/Jimmy_Osmond
Jimmy Page	http://en.wikipedia.org/wiki/Jimmy_Page
Jimmy Pop	http://en.wikipedia.org/wiki/Jimmy_Pop
Jimmy Smith	http://en.wikipedia.org/wiki/Jimmy_Smith_(musician)
Jimmy Smits	http://en.wikipedia.org/wiki/Jimmy_Smits
Jimmy Stewart	http://en.wikipedia.org/wiki/Jimmy_Stewart
Jimmy Swaggart	http://en.wikipedia.org/wiki/Jimmy_Swaggart
Jimmy The Greek	http://en.wikipedia.org/wiki/Jimmy_The_Greek
Jimmy Webb	http://en.wikipedia.org/wiki/Jimmy_Webb
Jiri Paroubek	http://en.wikipedia.org/wiki/Jiri_Paroubek
Jir� Paroubek	http://en.wikipedia.org/wiki/Jir%ED_Paroubek
Jo Ann Davis	http://en.wikipedia.org/wiki/Jo_Ann_Davis
Jo Ann Emerson	http://en.wikipedia.org/wiki/Jo_Ann_Emerson
Jo Anne Worley	http://en.wikipedia.org/wiki/Jo_Anne_Worley
Jo Bonner	http://en.wikipedia.org/wiki/Jo_Bonner
Jo Dee Messina	http://en.wikipedia.org/wiki/Jo_Dee_Messina
Jo Frost	http://en.wikipedia.org/wiki/Jo_Frost
Jo Johnson	http://en.wikipedia.org/wiki/Jo_Johnson
Jo Swinson	http://en.wikipedia.org/wiki/Jo_Swinson
Jo Van Fleet	http://en.wikipedia.org/wiki/Jo_Van_Fleet
Joachim du Bellay	http://en.wikipedia.org/wiki/Joachim_du_Bellay
Joachim von Ribbentrop	http://en.wikipedia.org/wiki/Joachim_von_Ribbentrop
Joan Allen	http://en.wikipedia.org/wiki/Joan_Allen
Joan Armatrading	http://en.wikipedia.org/wiki/Joan_Armatrading
Joan B. Kroc	http://en.wikipedia.org/wiki/Joan_B._Kroc
Joan Baez	http://en.wikipedia.org/wiki/Joan_Baez
Joan Baez	http://en.wikipedia.org/wiki/Joan_Baez
Joan Bennett	http://en.wikipedia.org/wiki/Joan_Bennett
Joan Blades	http://en.wikipedia.org/wiki/Joan_Blades
Joan Blondell	http://en.wikipedia.org/wiki/Joan_Blondell
Joan Caulfield	http://en.wikipedia.org/wiki/Joan_Caulfield
Joan Chen	http://en.wikipedia.org/wiki/Joan_Chen
Joan Collins	http://en.wikipedia.org/wiki/Joan_Collins
Joan Crawford	http://en.wikipedia.org/wiki/Joan_Crawford
Joan Cusack	http://en.wikipedia.org/wiki/Joan_Cusack
Joan D. Vinge	http://en.wikipedia.org/wiki/Joan_D._Vinge
Joan Davis	http://en.wikipedia.org/wiki/Joan_Davis
Joan Didion	http://en.wikipedia.org/wiki/Joan_Didion
Joan Enric Vives Sic�lia	http://en.wikipedia.org/wiki/Joan_Enric_Vives_Sic%EDlia
Joan Fontaine	http://en.wikipedia.org/wiki/Joan_Fontaine
Joan Gabriel Estany	http://en.wikipedia.org/wiki/Joan_Gabriel_i_Estany
Joan Ganz Cooney	http://en.wikipedia.org/wiki/Joan_Ganz_Cooney
Joan Hackett	http://en.wikipedia.org/wiki/Joan_Hackett
Joan Jett	http://en.wikipedia.org/wiki/Joan_Jett
Joan Kennedy	http://en.wikipedia.org/wiki/Joan_Kennedy
Joan Leslie	http://en.wikipedia.org/wiki/Joan_Leslie
Joan Lunden	http://en.wikipedia.org/wiki/Joan_Lunden
Joan Marsh	http://en.wikipedia.org/wiki/Joan_Marsh
Joan Mir�	http://en.wikipedia.org/wiki/Joan_Mir%F3
Joan of Arc	http://en.wikipedia.org/wiki/Joan_of_Arc
Joan Plowright	http://en.wikipedia.org/wiki/Joan_Plowright
Joan Rivers	http://en.wikipedia.org/wiki/Joan_Rivers
Joan Ruddock	http://en.wikipedia.org/wiki/Joan_Ruddock
Joan Severance	http://en.wikipedia.org/wiki/Joan_Severance
Joan Sutherland	http://en.wikipedia.org/wiki/Joan_Sutherland
Joan Van Ark	http://en.wikipedia.org/wiki/Joan_Van_Ark
Joan Walley	http://en.wikipedia.org/wiki/Joan_Walley
Joanna Baillie	http://en.wikipedia.org/wiki/Joanna_Baillie
Joanna Barnes	http://en.wikipedia.org/wiki/Joanna_Barnes
Joanna Cassidy	http://en.wikipedia.org/wiki/Joanna_Cassidy
Joanna Kerns	http://en.wikipedia.org/wiki/Joanna_Kerns
Joanna Lumley	http://en.wikipedia.org/wiki/Joanna_Lumley
Joanna Newsom	http://en.wikipedia.org/wiki/Joanna_Newsom
Joanna Russ	http://en.wikipedia.org/wiki/Joanna_Russ
Joanne Dru	http://en.wikipedia.org/wiki/Joanne_Dru
Joanne Woodward	http://en.wikipedia.org/wiki/Joanne_Woodward
J�annes Eidesgaard	http://en.wikipedia.org/wiki/J�annes_Eidesgaard
Jo�o Batista de Almeida Garrett	http://en.wikipedia.org/wiki/Almeida_Garrett
Jo�o Bernardo Vieira	http://en.wikipedia.org/wiki/Jo�o_Bernardo_Vieira
Jo�o de Deus	http://en.wikipedia.org/wiki/Jo�o_de_Deus
Jo�o I	http://en.wikipedia.org/wiki/John_I_of_Portugal
Jo�o II	http://en.wikipedia.org/wiki/John_II_of_Portugal
Jo�o III	http://en.wikipedia.org/wiki/John_III_of_Portugal
Jo�o IV	http://en.wikipedia.org/wiki/John_IV_of_Portugal
Jo�o V	http://en.wikipedia.org/wiki/John_V_of_Portugal
Jo�o VI	http://en.wikipedia.org/wiki/John_VI_of_Portugal
Joaquim Rafael Branco	http://en.wikipedia.org/wiki/Joaquim_Rafael_Branco
Joaquin Almunia	http://en.wikipedia.org/wiki/Joaquin_Almunia
Joaquin Miller	http://en.wikipedia.org/wiki/Joaquin_Miller
Joaquin Phoenix	http://en.wikipedia.org/wiki/Joaquin_Phoenix
JoBeth Williams	http://en.wikipedia.org/wiki/JoBeth_Williams
Jobyna Ralston	http://en.wikipedia.org/wiki/Jobyna_Ralston
Jock Mahoney	http://en.wikipedia.org/wiki/Jock_Mahoney
Jock Sturges	http://en.wikipedia.org/wiki/Jock_Sturges
Jodi Lyn O'Keefe	http://en.wikipedia.org/wiki/Jodi_Lyn_O%27Keefe
Jodi Rell	http://en.wikipedia.org/wiki/Jodi_Rell
Jodie Foster	http://en.wikipedia.org/wiki/Jodie_Foster
Jodie Marsh	http://en.wikipedia.org/wiki/Jodie_Marsh
Jodie Sweetin	http://en.wikipedia.org/wiki/Jodie_Sweetin
Jody Miller	http://en.wikipedia.org/wiki/Jody_Miller
Jody Powell	http://en.wikipedia.org/wiki/Jody_Powell
Jody Watley	http://en.wikipedia.org/wiki/Jody_Watley
Jody Williams	http://en.wikipedia.org/wiki/Jody_Williams
Joe Absolom	http://en.wikipedia.org/wiki/Joe_Absolom
Joe Adonis	http://en.wikipedia.org/wiki/Joe_Adonis
Joe Allbaugh	http://en.wikipedia.org/wiki/Joe_Allbaugh
Joe Allison	http://en.wikipedia.org/wiki/Joe_Allison
Joe Arpaio	http://en.wikipedia.org/wiki/Joe_Arpaio
Joe Baca	http://en.wikipedia.org/wiki/Joe_Baca
Joe Barton	http://en.wikipedia.org/wiki/Joe_Barton
Joe Barton	http://en.wikipedia.org/wiki/Joe_Barton
Joe Benton	http://en.wikipedia.org/wiki/Joe_Benton
Joe Besser	http://en.wikipedia.org/wiki/Joe_Besser
Joe Bob Briggs	http://en.wikipedia.org/wiki/Joe_Bob_Briggs
Joe Budden	http://en.wikipedia.org/wiki/Joe_Budden
Joe C.	http://en.wikipedia.org/wiki/Joe_C.
Joe Clark	http://en.wikipedia.org/wiki/Joe_Clark
Joe Cocker	http://en.wikipedia.org/wiki/Joe_Cocker
Joe Conason	http://en.wikipedia.org/wiki/Joe_Conason
Joe Coulombe	http://en.wikipedia.org/wiki/Joe_Coulombe
Joe Courtney	http://en.wikipedia.org/wiki/Joe_Courtney_(politician)
Joe Cronin	http://en.wikipedia.org/wiki/Joe_Cronin
Joe Dallesandro	http://en.wikipedia.org/wiki/Joe_Dallesandro
Joe Dante	http://en.wikipedia.org/wiki/Joe_Dante
Joe DeRita	http://en.wikipedia.org/wiki/Joe_DeRita
Joe DiMaggio	http://en.wikipedia.org/wiki/Joe_DiMaggio
Joe Don Baker	http://en.wikipedia.org/wiki/Joe_Don_Baker
Joe Donnelly	http://en.wikipedia.org/wiki/Joe_Donnelly
Joe E. Brown	http://en.wikipedia.org/wiki/Joe_E._Brown_(comedian)
Joe E. Ross	http://en.wikipedia.org/wiki/Joe_E._Ross
Joe Elliott	http://en.wikipedia.org/wiki/Joe_Elliott
Joe Eszterhas	http://en.wikipedia.org/wiki/Joe_Eszterhas
Joe Flaherty	http://en.wikipedia.org/wiki/Joe_Flaherty
Joe Flanigan	http://en.wikipedia.org/wiki/Joe_Flanigan
Joe Francis	http://en.wikipedia.org/wiki/Joe_Francis
Joe Franklin	http://en.wikipedia.org/wiki/Joe_Franklin
Joe Frazier	http://en.wikipedia.org/wiki/Joe_Frazier
Joe Garagiola	http://en.wikipedia.org/wiki/Joe_Garagiola
Joe Gold	http://en.wikipedia.org/wiki/Joe_Gold
Joe Hill	http://en.wikipedia.org/wiki/Joe_Hill
Joe Jackson	http://en.wikipedia.org/wiki/Joe_Jackson_(musician)
Joe Jackson	http://en.wikipedia.org/wiki/Joe_Jackson_(manager)
Joe Johnston	http://en.wikipedia.org/wiki/Joe_Johnston
Joe Klein	http://en.wikipedia.org/wiki/Joe_Klein
Joe Kolter	http://en.wikipedia.org/wiki/Joe_Kolter
Joe Lando	http://en.wikipedia.org/wiki/Joe_Lando
Joe Lo Truglio	http://en.wikipedia.org/wiki/Joe_Lo_Truglio
Joe Lockhart	http://en.wikipedia.org/wiki/Joe_Lockhart
Joe Louis	http://en.wikipedia.org/wiki/Joe_Louis
Joe Manchin	http://en.wikipedia.org/wiki/Joe_Manchin
Joe Mantegna	http://en.wikipedia.org/wiki/Joe_Mantegna
Joe Masseria	http://en.wikipedia.org/wiki/Joe_Masseria
Joe McCarthy	http://en.wikipedia.org/wiki/Joe_McCarthy_(manager)
Joe Meek	http://en.wikipedia.org/wiki/Joe_Meek
Joe Montana	http://en.wikipedia.org/wiki/Joe_Montana
Joe Morgan	http://en.wikipedia.org/wiki/Joe_Morgan
Joe Morton	http://en.wikipedia.org/wiki/Joe_Morton
Joe Namath	http://en.wikipedia.org/wiki/Joe_Namath
Joe Orton	http://en.wikipedia.org/wiki/Joe_Orton
Joe Pantoliano	http://en.wikipedia.org/wiki/Joe_Pantoliano
Joe Paterno	http://en.wikipedia.org/wiki/Joe_Paterno
Joe Penner	http://en.wikipedia.org/wiki/Joe_Penner
Joe Penny	http://en.wikipedia.org/wiki/Joe_Penny
Joe Perry	http://en.wikipedia.org/wiki/Joe_Perry_(musician)
Joe Pesci	http://en.wikipedia.org/wiki/Joe_Pesci
Joe Piscopo	http://en.wikipedia.org/wiki/Joe_Piscopo
Joe Regalbuto	http://en.wikipedia.org/wiki/Joe_Regalbuto
Joe Rogan	http://en.wikipedia.org/wiki/Joe_Rogan
Joe Roth	http://en.wikipedia.org/wiki/Joe_Roth
Joe Sacco	http://en.wikipedia.org/wiki/Joe_Sacco
Joe Santos	http://en.wikipedia.org/wiki/Joe_Santos
Joe Satriani	http://en.wikipedia.org/wiki/Joe_Satriani
Joe Sawyer	http://en.wikipedia.org/wiki/Joe_Sawyer
Joe Scarborough	http://en.wikipedia.org/wiki/Joe_Scarborough
Joe Schermie	http://en.wikipedia.org/wiki/Joe_Schermie
Joe Schwarz	http://en.wikipedia.org/wiki/Joe_Schwarz
Joe Sestak	http://en.wikipedia.org/wiki/Joe_Sestak
Joe Skeen	http://en.wikipedia.org/wiki/Joe_Skeen
Joe Spano	http://en.wikipedia.org/wiki/Joe_Spano
Joe Spinell	http://en.wikipedia.org/wiki/Joe_Spinell
Joe Strummer	http://en.wikipedia.org/wiki/Joe_Strummer
Joe Theismann	http://en.wikipedia.org/wiki/Joe_Theismann
Joe Torre	http://en.wikipedia.org/wiki/Joe_Torre
Joe Viterelli	http://en.wikipedia.org/wiki/Joe_Viterelli
Joe Walsh	http://en.wikipedia.org/wiki/Joe_Walsh
Joe Wilson	http://en.wikipedia.org/wiki/Joe_Wilson_(U.S._politician)
Joel Barlow	http://en.wikipedia.org/wiki/Joel_Barlow
Joel Chandler Harris	http://en.wikipedia.org/wiki/Joel_Chandler_Harris
Joel Coen	http://en.wikipedia.org/wiki/Joel_Coen
Joel D. Kaplan	http://en.wikipedia.org/wiki/Joel_Kaplan
Joel Dorius	http://en.wikipedia.org/wiki/Joel_Dorius
Joel Elias Spingarn	http://en.wikipedia.org/wiki/Joel_Elias_Spingarn
Joel Gretsch	http://en.wikipedia.org/wiki/Joel_Gretsch
Joel Grey	http://en.wikipedia.org/wiki/Joel_Grey
Joel Hefley	http://en.wikipedia.org/wiki/Joel_Hefley
Joel Hodgson	http://en.wikipedia.org/wiki/Joel_Hodgson
Joel Madden	http://en.wikipedia.org/wiki/Joel_Madden
Joel McCrea	http://en.wikipedia.org/wiki/Joel_McCrea
Joel Schumacher	http://en.wikipedia.org/wiki/Joel_Schumacher
Joel Siegel	http://en.wikipedia.org/wiki/Joel_Siegel
Joel-Peter Witkin	http://en.wikipedia.org/wiki/Joel-Peter_Witkin
Joely Fisher	http://en.wikipedia.org/wiki/Joely_Fisher
Joely Richardson	http://en.wikipedia.org/wiki/Joely_Richardson
Joergen Nash	http://en.wikipedia.org/wiki/Joergen_Nash
Joey Bishop	http://en.wikipedia.org/wiki/Joey_Bishop
Joey Buttafuoco	http://en.wikipedia.org/wiki/Joey_Buttafuoco
Joey Fatone	http://en.wikipedia.org/wiki/Joey_Fatone
Joey Heatherton	http://en.wikipedia.org/wiki/Joey_Heatherton
Joey Jordison	http://en.wikipedia.org/wiki/Joey_Jordison
Joey Lauren Adams	http://en.wikipedia.org/wiki/Joey_Lauren_Adams
Joey Lawrence	http://en.wikipedia.org/wiki/Joey_Lawrence
Joey McIntyre	http://en.wikipedia.org/wiki/Joey_McIntyre
Joey Ramone	http://en.wikipedia.org/wiki/Joey_Ramone
Joey Santiago	http://en.wikipedia.org/wiki/Joey_Santiago
Joey Skaggs	http://en.wikipedia.org/wiki/Joey_Skaggs
Joh Bjelke-Petersen	http://en.wikipedia.org/wiki/Joh_Bjelke-Petersen
Johan Cruijff	http://en.wikipedia.org/wiki/Johan_Cruijff
Johan de Witt	http://en.wikipedia.org/wiki/Johan_de_Witt
Johan Helsingius	http://en.wikipedia.org/wiki/Johan_Helsingius
Johan Sverdrup	http://en.wikipedia.org/wiki/Johan_Sverdrup
Johann Adolph Hasse	http://en.wikipedia.org/wiki/Johann_Adolph_Hasse
Johann Augustus Eberhard	http://en.wikipedia.org/wiki/Johann_Augustus_Eberhard
Johann Baptist Cramer	http://en.wikipedia.org/wiki/Johann_Baptist_Cramer
Johann Christian Fabricius	http://en.wikipedia.org/wiki/Johann_Christian_Fabricius
Johann Christian Poggendorff	http://en.wikipedia.org/wiki/Johann_Christian_Poggendorff
Johann Deisenhofer	http://en.wikipedia.org/wiki/Johann_Deisenhofer
Johann Eck	http://en.wikipedia.org/wiki/Johann_Eck
Johann Franz Encke	http://en.wikipedia.org/wiki/Johann_Franz_Encke
Johann Friedrich Overbeck	http://en.wikipedia.org/wiki/Johann_Friedrich_Overbeck
Johann Friedrich Struensee	http://en.wikipedia.org/wiki/Johann_Friedrich_Struensee
Johann Georg Hamann	http://en.wikipedia.org/wiki/Johann_Georg_Hamann
Johann Gottfried Eichhorn	http://en.wikipedia.org/wiki/Johann_Gottfried_Eichhorn
Johann Gottfried Herder	http://en.wikipedia.org/wiki/Johann_Gottfried_Herder
Johann Gottlieb Fichte	http://en.wikipedia.org/wiki/Johann_Gottlieb_Fichte
Johann Heinrich Lambert	http://en.wikipedia.org/wiki/Johann_Heinrich_Lambert
Johann Heinrich Pestalozzi	http://en.wikipedia.org/wiki/Johann_Heinrich_Pestalozzi
Johann Jakob Bodmer	http://en.wikipedia.org/wiki/Johann_Jakob_Bodmer
Johann Joseph Fux	http://en.wikipedia.org/wiki/Johann_Joseph_Fux
Johann Kaspar Lavater	http://en.wikipedia.org/wiki/Johann_Kaspar_Lavater
Johann Nikolaus von Hontheim	http://en.wikipedia.org/wiki/Johann_Nikolaus_von_Hontheim
Johann Pachelbel	http://en.wikipedia.org/wiki/Johann_Pachelbel
Johann Reuchlin	http://en.wikipedia.org/wiki/Johann_Reuchlin
Johann Sebastian Bach	http://en.wikipedia.org/wiki/Johann_Sebastian_Bach
Johann Strauss	http://en.wikipedia.org/wiki/Johann_Strauss_II
Johann Strauss, Sr.	http://en.wikipedia.org/wiki/Johann_Strauss%2C_Sr.
Johann Tauler	http://en.wikipedia.org/wiki/Johann_Tauler
Johann Tetzel	http://en.wikipedia.org/wiki/Johann_Tetzel
Johann Tobias Mayer	http://en.wikipedia.org/wiki/Tobias_Mayer
Johann Winckelmann	http://en.wikipedia.org/wiki/Johann_Winckelmann
J�hanna Sigur�ard�ttir	http://en.wikipedia.org/wiki/J�hanna_Sigur�ard�ttir
Johannes Brahms	http://en.wikipedia.org/wiki/Johannes_Brahms
Johannes Carsten Hauch	http://en.wikipedia.org/wiki/Johannes_Carsten_Hauch
Johannes Diderik van der Waals	http://en.wikipedia.org/wiki/Johannes_Diderik_van_der_Waals
Johannes Gutenberg	http://en.wikipedia.org/wiki/Johannes_Gutenberg
Johannes Heesters	http://en.wikipedia.org/wiki/Johannes_Heesters
Johannes Hevelius	http://en.wikipedia.org/wiki/Johannes_Hevelius
Johannes Kepler	http://en.wikipedia.org/wiki/Johannes_Kepler
Johannes Popitz	http://en.wikipedia.org/wiki/Johannes_Popitz
Johannes Rau	http://en.wikipedia.org/wiki/Johannes_Rau
Johannes Rydberg	http://en.wikipedia.org/wiki/Johannes_Rydberg
Johannes Scotus Erigena	http://en.wikipedia.org/wiki/Johannes_Scotus_Erigena
Johannes Stark	http://en.wikipedia.org/wiki/Johannes_Stark
Johannes Stumpf	http://en.wikipedia.org/wiki/Johann_Stumpf_(writer)
Johannes Wier	http://en.wikipedia.org/wiki/Johannes_Wier
John 5	http://en.wikipedia.org/wiki/John_5_(guitarist)
John A. Luke Jr.	http://en.wikipedia.org/wiki/John_A._Luke_Jr.
John A. Macdonald	http://en.wikipedia.org/wiki/John_A._Macdonald
John A. Pople	http://en.wikipedia.org/wiki/John_A._Pople
John A. Quitman	http://en.wikipedia.org/wiki/John_A._Quitman
John Abbott	http://en.wikipedia.org/wiki/John_Abbott
John Abizaid	http://en.wikipedia.org/wiki/John_Abizaid
John Abraham	http://en.wikipedia.org/wiki/John_Abraham_(actor)
John Adams	http://en.wikipedia.org/wiki/John_Adams
John Adams Dix	http://en.wikipedia.org/wiki/John_Adams_Dix
John Addington Symonds	http://en.wikipedia.org/wiki/John_Addington_Symonds
John Addison	http://en.wikipedia.org/wiki/John_Addison
John Adler	http://en.wikipedia.org/wiki/John_Adler
John Agar	http://en.wikipedia.org/wiki/John_Agar
John Albert Carroll	http://en.wikipedia.org/wiki/John_Albert_Carroll
John Ales	http://en.wikipedia.org/wiki/John_Ales
John Alexander	http://en.wikipedia.org/wiki/John_Alexander_(actor)
John Alexander McClernand	http://en.wikipedia.org/wiki/John_Alexander_McClernand
John Alexander Reina Newlands	http://en.wikipedia.org/wiki/John_Alexander_Reina_Newlands
John Alford	http://en.wikipedia.org/wiki/John_Alford_(actor)
John Allen Muhammad	http://en.wikipedia.org/wiki/John_Allen_Muhammad
John Altman	http://en.wikipedia.org/wiki/John_Altman_(actor)
John Amos	http://en.wikipedia.org/wiki/John_Amos
John Anderson	http://en.wikipedia.org/wiki/John_Anderson_(musician)
John Anderson	http://en.wikipedia.org/wiki/John_B._Anderson
John Aniston	http://en.wikipedia.org/wiki/John_Aniston
John Ankerberg	http://en.wikipedia.org/wiki/John_Ankerberg
John Aprea	http://en.wikipedia.org/wiki/John_Aprea
John Arbuthnot	http://en.wikipedia.org/wiki/John_Arbuthnot
John Archibald Wheeler	http://en.wikipedia.org/wiki/John_Archibald_Wheeler
John Arden	http://en.wikipedia.org/wiki/John_Arden
John Armstrong	http://en.wikipedia.org/wiki/John_Armstrong,_Jr.
John Ashbery	http://en.wikipedia.org/wiki/John_Ashbery
John Ashcroft	http://en.wikipedia.org/wiki/John_Ashcroft
John Astin	http://en.wikipedia.org/wiki/John_Astin
John Atta Mills	http://en.wikipedia.org/wiki/John_Atta_Mills
John B. Breaux	http://en.wikipedia.org/wiki/John_B._Breaux
John B. Fenn	http://en.wikipedia.org/wiki/John_B._Fenn
John B. Hess	http://en.wikipedia.org/wiki/John_B._Hess
John Bach McMaster	http://en.wikipedia.org/wiki/John_Bach_McMaster
John Badham	http://en.wikipedia.org/wiki/John_Badham
John Bainbridge	http://en.wikipedia.org/wiki/John_Bainbridge_(astronomer)
John Balance	http://en.wikipedia.org/wiki/John_Balance
John Baldacci	http://en.wikipedia.org/wiki/John_Baldacci
John Baldacci	http://en.wikipedia.org/wiki/John_Baldacci
John Ball	http://en.wikipedia.org/wiki/John_Ball_(priest)
John Ball	http://en.wikipedia.org/wiki/John_Ball_(naturalist)
John Banner	http://en.wikipedia.org/wiki/John_Banner
John Banville	http://en.wikipedia.org/wiki/John_Banville
John Bardeen	http://en.wikipedia.org/wiki/John_Bardeen
John Baron	http://en.wikipedia.org/wiki/John_Baron_(MP)
John Barrasso	http://en.wikipedia.org/wiki/John_Barrasso
John Barrow	http://en.wikipedia.org/wiki/John_Barrow_(U.S._politician)
John Barrowman	http://en.wikipedia.org/wiki/John_Barrowman
John Barry	http://en.wikipedia.org/wiki/John_Barry_(composer)
John Barrymore	http://en.wikipedia.org/wiki/John_Barrymore
John Barth	http://en.wikipedia.org/wiki/John_Barth
John Bartlett	http://en.wikipedia.org/wiki/John_Bartlett_(publisher)
John Bates Clark	http://en.wikipedia.org/wiki/John_Bates_Clark
John Battelle	http://en.wikipedia.org/wiki/John_Battelle
John Bayley	http://en.wikipedia.org/wiki/John_Bayley_(writer)
John Beal	http://en.wikipedia.org/wiki/John_Beal_(actor)
John Bell Hood	http://en.wikipedia.org/wiki/John_Bell_Hood
John Belushi	http://en.wikipedia.org/wiki/John_Belushi
John Bercow	http://en.wikipedia.org/wiki/John_Bercow
John Berger	http://en.wikipedia.org/wiki/John_Berger
John Bernard Burke	http://en.wikipedia.org/wiki/John_Bernard_Burke
John Berryman	http://en.wikipedia.org/wiki/John_Berryman
John Betjeman	http://en.wikipedia.org/wiki/John_Betjeman
John Biddle	http://en.wikipedia.org/wiki/John_Biddle_(Unitarian)
John Bigelow	http://en.wikipedia.org/wiki/John_Bigelow
John Birch	http://en.wikipedia.org/wiki/John_Birch_(missionary)
John Blow	http://en.wikipedia.org/wiki/John_Blow
John Boccieri	http://en.wikipedia.org/wiki/John_Boccieri
John Boehner	http://en.wikipedia.org/wiki/John_Boehner
John Bolton	http://en.wikipedia.org/wiki/John_R._Bolton
John Bonham	http://en.wikipedia.org/wiki/John_Bonham
John Boorman	http://en.wikipedia.org/wiki/John_Boorman
John Boozman	http://en.wikipedia.org/wiki/John_Boozman
John Bowen	http://en.wikipedia.org/wiki/John_Griffith_Bowen
John Boyd Orr	http://en.wikipedia.org/wiki/John_Boyd_Orr
John Brademas	http://en.wikipedia.org/wiki/John_Brademas
John Bradshaw	http://en.wikipedia.org/wiki/John_Bradshaw_(judge)
John Braine	http://en.wikipedia.org/wiki/John_Braine
John Brand	http://en.wikipedia.org/wiki/John_Brand
John Breaux	http://en.wikipedia.org/wiki/John_Breaux
John Brockington	http://en.wikipedia.org/wiki/John_Brockington
John Brockman	http://en.wikipedia.org/wiki/John_Brockman_(literary_agent)
John Brogden	http://en.wikipedia.org/wiki/John_Brogden_(politician)
John Bromfield	http://en.wikipedia.org/wiki/John_Bromfield
John Brougham	http://en.wikipedia.org/wiki/John_Brougham
John Brown	http://en.wikipedia.org/wiki/John_Brown_(abolitionist)
John Browne	http://en.wikipedia.org/wiki/John_Browne,_Baron_Browne_of_Madingley
John Browning	http://en.wikipedia.org/wiki/John_Browning
John Brunner	http://en.wikipedia.org/wiki/John_Brunner_(novelist)
John Bruton	http://en.wikipedia.org/wiki/John_Bruton
John Bryan	http://en.wikipedia.org/wiki/John_Bryan_(diplomat)
John Bryant	http://en.wikipedia.org/wiki/John_Wiley_Bryant
John Buchan	http://en.wikipedia.org/wiki/John_Buchan
John Bull	http://en.wikipedia.org/wiki/John_Bull_(composer)
John Bunnell	http://en.wikipedia.org/wiki/John_Bunnell
John Bunny	http://en.wikipedia.org/wiki/John_Bunny
John Bunyan	http://en.wikipedia.org/wiki/John_Bunyan
John Burgoyne	http://en.wikipedia.org/wiki/John_Burgoyne
John Burns	http://en.wikipedia.org/wiki/John_F._Burns
John Burroughs	http://en.wikipedia.org/wiki/John_Burroughs
John Byner	http://en.wikipedia.org/wiki/John_Byner
John C. Breckinridge	http://en.wikipedia.org/wiki/John_C._Breckinridge
John C. Calhoun	http://en.wikipedia.org/wiki/John_C._Calhoun
John C. Danforth	http://en.wikipedia.org/wiki/John_C._Danforth
John C. Fleming	http://en.wikipedia.org/wiki/John_C._Fleming
John C. Fremont	http://en.wikipedia.org/wiki/John_C._Fremont
John C. Kendrew	http://en.wikipedia.org/wiki/John_C._Kendrew
John C. Polanyi	http://en.wikipedia.org/wiki/John_C._Polanyi
John C. Reilly	http://en.wikipedia.org/wiki/John_C._Reilly
John C. Stennis	http://en.wikipedia.org/wiki/John_C._Stennis
John C. Whitehead	http://en.wikipedia.org/wiki/John_C._Whitehead
John Cabot	http://en.wikipedia.org/wiki/John_Cabot
John Cage	http://en.wikipedia.org/wiki/John_Cage
John Caius	http://en.wikipedia.org/wiki/John_Caius
John Cale	http://en.wikipedia.org/wiki/John_Cale
John Callcott Horsley	http://en.wikipedia.org/wiki/John_Callcott_Horsley
John Calvin	http://en.wikipedia.org/wiki/John_Calvin
John Cameron	http://en.wikipedia.org/wiki/John_Cameron_(theologian)
John Cameron Mitchell	http://en.wikipedia.org/wiki/John_Cameron_Mitchell
John Campbell	http://en.wikipedia.org/wiki/John_B._T._Campbell_III
John Candy	http://en.wikipedia.org/wiki/John_Candy
John Cardinal O'Connor	http://en.wikipedia.org/wiki/John_Cardinal_O%27Connor
John Carmack	http://en.wikipedia.org/wiki/John_Carmack
John Carpenter	http://en.wikipedia.org/wiki/John_Carpenter
John Carradine	http://en.wikipedia.org/wiki/John_Carradine
John Carter	http://en.wikipedia.org/wiki/John_Carter_(Texas)
John Cassavetes	http://en.wikipedia.org/wiki/John_Cassavetes
John Cassell	http://en.wikipedia.org/wiki/John_Cassell
John Cavanaugh	http://en.wikipedia.org/wiki/John_Joseph_Cavanaugh_III
John Cazale	http://en.wikipedia.org/wiki/John_Cazale
John Cena	http://en.wikipedia.org/wiki/John_Cena
John Chancellor	http://en.wikipedia.org/wiki/John_Chancellor
John Charles Daly	http://en.wikipedia.org/wiki/John_Charles_Daly
John Cheever	http://en.wikipedia.org/wiki/John_Cheever
John Cho	http://en.wikipedia.org/wiki/John_Cho
John Ciardi	http://en.wikipedia.org/wiki/John_Ciardi
John Clare	http://en.wikipedia.org/wiki/John_Clare
John Cleese	http://en.wikipedia.org/wiki/John_Cleese
John Cockcroft	http://en.wikipedia.org/wiki/John_Cockcroft
John Coltrane	http://en.wikipedia.org/wiki/John_Coltrane
John Connally	http://en.wikipedia.org/wiki/John_Connally
John Constable	http://en.wikipedia.org/wiki/John_Constable
John Conway	http://en.wikipedia.org/wiki/John_Horton_Conway
John Conyers	http://en.wikipedia.org/wiki/John_Conyers
John Conyers, Jr.	http://en.wikipedia.org/wiki/John_Conyers%2C_Jr.
John Corbett	http://en.wikipedia.org/wiki/John_Corbett_(actor)
John Cornforth	http://en.wikipedia.org/wiki/John_Cornforth
John Cornyn	http://en.wikipedia.org/wiki/John_Cornyn
John Costello	http://en.wikipedia.org/wiki/John_Costello
John Cotton	http://en.wikipedia.org/wiki/John_Cotton_(Puritan)
John Couch Adams	http://en.wikipedia.org/wiki/John_Couch_Adams
John Cougar Mellencamp	http://en.wikipedia.org/wiki/John_Cougar_Mellencamp
John Cowper Powys	http://en.wikipedia.org/wiki/John_Cowper_Powys
John Crome	http://en.wikipedia.org/wiki/John_Crome
John Cromwell	http://en.wikipedia.org/wiki/John_Cromwell_(director)
John Crowe Ransom	http://en.wikipedia.org/wiki/John_Crowe_Ransom
John Cryer	http://en.wikipedia.org/wiki/John_Cryer
John Culberson	http://en.wikipedia.org/wiki/John_Culberson
John Cullum	http://en.wikipedia.org/wiki/John_Cullum
John Cusack	http://en.wikipedia.org/wiki/John_Cusack
John D. Dingell	http://en.wikipedia.org/wiki/John_D._Dingell
John D. MacArthur	http://en.wikipedia.org/wiki/John_D._MacArthur
John D. MacDonald	http://en.wikipedia.org/wiki/John_D._MacDonald
John D. Roberts	http://en.wikipedia.org/wiki/John_Roberts_(television_reporter)
John D. Rockefeller	http://en.wikipedia.org/wiki/John_D._Rockefeller
John D. Rockefeller IV	http://en.wikipedia.org/wiki/John_D._Rockefeller_IV
John D. Rockefeller, Jr.	http://en.wikipedia.org/wiki/John_D._Rockefeller%2C_Jr.
John Dalton	http://en.wikipedia.org/wiki/John_Dalton
John Daly	http://en.wikipedia.org/wiki/John_Daly_(golfer)
John Danforth	http://en.wikipedia.org/wiki/John_Danforth
John Davidson	http://en.wikipedia.org/wiki/John_Davidson_(entertainer)
John Davis	http://en.wikipedia.org/wiki/John_Davis_(English_explorer)
John Day	http://en.wikipedia.org/wiki/John_Day_(dramatist)
John de Stratford	http://en.wikipedia.org/wiki/John_de_Stratford
John Deacon	http://en.wikipedia.org/wiki/John_Deacon
John Dean	http://en.wikipedia.org/wiki/John_Dean
John Dee	http://en.wikipedia.org/wiki/John_Dee
John DeLorean	http://en.wikipedia.org/wiki/John_DeLorean
John Demjanjuk	http://en.wikipedia.org/wiki/John_Demjanjuk
John Denham	http://en.wikipedia.org/wiki/John_Denham_(politician)
John Dennis	http://en.wikipedia.org/wiki/John_Dennis_(dramatist)
John Densmore	http://en.wikipedia.org/wiki/John_Densmore
John Denver	http://en.wikipedia.org/wiki/John_Denver
John Derek	http://en.wikipedia.org/wiki/John_Derek
John Deutch	http://en.wikipedia.org/wiki/John_Deutch
John Dewey	http://en.wikipedia.org/wiki/John_Dewey
John Dickerson	http://en.wikipedia.org/wiki/John_Dickerson_(journalist)
John Dickinson	http://en.wikipedia.org/wiki/John_Dickinson_(delegate)
John Diebold	http://en.wikipedia.org/wiki/John_Diebold
John Diefenbaker	http://en.wikipedia.org/wiki/John_Diefenbaker
John Diehl	http://en.wikipedia.org/wiki/John_Diehl
John Dillinger	http://en.wikipedia.org/wiki/John_Dillinger
John Dingell	http://en.wikipedia.org/wiki/John_Dingell
John Doe	http://en.wikipedia.org/wiki/John_Doe_(musician)
John Doerr	http://en.wikipedia.org/wiki/John_Doerr
John Dollond	http://en.wikipedia.org/wiki/John_Dollond
John Doman	http://en.wikipedia.org/wiki/John_Doman
John Donne	http://en.wikipedia.org/wiki/John_Donne
John Doolittle	http://en.wikipedia.org/wiki/John_Doolittle
John Dos Passos	http://en.wikipedia.org/wiki/John_Dos_Passos
John Dowland	http://en.wikipedia.org/wiki/John_Dowland
John Drew Barrymore	http://en.wikipedia.org/wiki/John_Drew_Barrymore
John Dryden	http://en.wikipedia.org/wiki/John_Dryden
John Duncan	http://en.wikipedia.org/wiki/Jimmy_Duncan_(U.S._politician)
John Duns Scotus	http://en.wikipedia.org/wiki/John_Duns_Scotus
John Dvorak	http://en.wikipedia.org/wiki/John_Dvorak
John Dye	http://en.wikipedia.org/wiki/John_Dye
John E. du Pont	http://en.wikipedia.org/wiki/John_E._du_Pont
John E. Grotberg	http://en.wikipedia.org/wiki/John_E._Grotberg
John E. McLaughlin	http://en.wikipedia.org/wiki/John_E._McLaughlin
John E. O'Neill	http://en.wikipedia.org/wiki/John_E._O%27Neill
John E. Sununu	http://en.wikipedia.org/wiki/John_E._Sununu
John E. Walker	http://en.wikipedia.org/wiki/John_E._Walker
John Earle	http://en.wikipedia.org/wiki/John_Earle_(bishop)
John Edgar Wideman	http://en.wikipedia.org/wiki/John_Edgar_Wideman
John Edward	http://en.wikipedia.org/wiki/John_Edward
John Edward Porter	http://en.wikipedia.org/wiki/John_Edward_Porter
John Edward Robinson	http://en.wikipedia.org/wiki/John_Edward_Robinson_(serial_killer)
John Edwards	http://en.wikipedia.org/wiki/John_Edwards
John Ehrlichman	http://en.wikipedia.org/wiki/John_Ehrlichman
John Elway	http://en.wikipedia.org/wiki/John_Elway
John Engler	http://en.wikipedia.org/wiki/John_Engler
John Ennis	http://en.wikipedia.org/wiki/John_Ennis_(actor)
John Enos III	http://en.wikipedia.org/wiki/John_Enos_III
John Ensign	http://en.wikipedia.org/wiki/John_Ensign
John Entwistle	http://en.wikipedia.org/wiki/John_Entwistle
John Ericsson	http://en.wikipedia.org/wiki/John_Ericsson
John Erlenborn	http://en.wikipedia.org/wiki/John_Erlenborn
John Evander Couey	http://en.wikipedia.org/wiki/John_Evander_Couey
John Evelyn	http://en.wikipedia.org/wiki/John_Evelyn
John Everett Millais	http://en.wikipedia.org/wiki/John_Everett_Millais
John F. Akers	http://en.wikipedia.org/wiki/John_F._Akers
John F. Gifford	http://en.wikipedia.org/wiki/Jack_Gifford_(businessman)
John F. Kennedy	http://en.wikipedia.org/wiki/John_F._Kennedy
John F. Kennedy, Jr.	http://en.wikipedia.org/wiki/John_F._Kennedy%2C_Jr.
John F. Kerry	http://en.wikipedia.org/wiki/John_F._Kerry
John F. Lehman	http://en.wikipedia.org/wiki/John_F._Lehman
John F. Seiberling	http://en.wikipedia.org/wiki/John_F._Seiberling
John F. Street	http://en.wikipedia.org/wiki/John_F._Street
John Fahey	http://en.wikipedia.org/wiki/John_M._Fahey,_Jr.
John Fahey	http://en.wikipedia.org/wiki/John_Fahey_(musician)
John Fante	http://en.wikipedia.org/wiki/John_Fante
John Farrow	http://en.wikipedia.org/wiki/John_Farrow
John Fiedler	http://en.wikipedia.org/wiki/John_Fiedler
John Field	http://en.wikipedia.org/wiki/John_Field_(composer)
John Fiske	http://en.wikipedia.org/wiki/John_Fiske_(philosopher)
John Flamsteed	http://en.wikipedia.org/wiki/John_Flamsteed
John Flansburgh	http://en.wikipedia.org/wiki/John_Flansburgh
John Fogerty	http://en.wikipedia.org/wiki/John_Fogerty
John Ford	http://en.wikipedia.org/wiki/John_Ford
John Forster	http://en.wikipedia.org/wiki/John_Forster_(biographer)
John Forsythe	http://en.wikipedia.org/wiki/John_Forsythe
John Foster Dulles	http://en.wikipedia.org/wiki/John_Foster_Dulles
John Fowles	http://en.wikipedia.org/wiki/John_Fowles
John Foxe	http://en.wikipedia.org/wiki/John_Foxe
John Francis Lewis	http://en.wikipedia.org/wiki/John_Francis_Lewis
John Frankenheimer	http://en.wikipedia.org/wiki/John_Frankenheimer
John Freind	http://en.wikipedia.org/wiki/John_Freind
John Frusciante	http://en.wikipedia.org/wiki/John_Frusciante
John Fund	http://en.wikipedia.org/wiki/John_Fund
John G. Avildsen	http://en.wikipedia.org/wiki/John_G._Avildsen
John G. Brady	http://en.wikipedia.org/wiki/John_G._Brady
John G. Drosdick	http://en.wikipedia.org/wiki/John_Drosdick
John G. Neihardt	http://en.wikipedia.org/wiki/John_G._Neihardt
John G. Roberts, Jr.	http://en.wikipedia.org/wiki/John_G._Roberts%2C_Jr.
John G. Rowland	http://en.wikipedia.org/wiki/John_G._Rowland
John G. Schmitz	http://en.wikipedia.org/wiki/John_G._Schmitz
John Galliano	http://en.wikipedia.org/wiki/John_Galliano
John Galsworthy	http://en.wikipedia.org/wiki/John_Galsworthy
John Galt	http://en.wikipedia.org/wiki/John_Galt_(novelist)
John Garamendi	http://en.wikipedia.org/wiki/John_Garamendi
John Gardner	http://en.wikipedia.org/wiki/John_Gardner_(novelist)
John Garfield	http://en.wikipedia.org/wiki/John_Garfield
John Gavin	http://en.wikipedia.org/wiki/John_Gavin
John Gay	http://en.wikipedia.org/wiki/John_Gay
John Gibson	http://en.wikipedia.org/wiki/John_Gibson_(political_commentator)
John Gibson	http://en.wikipedia.org/wiki/John_Gibson_(sculptor)
John Gielgud	http://en.wikipedia.org/wiki/John_Gielgud
John Gilbert	http://en.wikipedia.org/wiki/John_Gilbert_(actor)
John Gilmore	http://en.wikipedia.org/wiki/John_Gilmore_(activist)
John Glen	http://en.wikipedia.org/wiki/John_Glen_(MP)
John Glenn	http://en.wikipedia.org/wiki/John_Glenn
John Glover	http://en.wikipedia.org/wiki/John_Glover_(actor)
John Goodman	http://en.wikipedia.org/wiki/John_Goodman
John Gotti	http://en.wikipedia.org/wiki/John_Gotti
John Greenleaf Whittier	http://en.wikipedia.org/wiki/John_Greenleaf_Whittier
John Gregory Dunne	http://en.wikipedia.org/wiki/John_Gregory_Dunne
John Gregson	http://en.wikipedia.org/wiki/John_Gregson
John Grisham	http://en.wikipedia.org/wiki/John_Grisham
John Guare	http://en.wikipedia.org/wiki/John_Guare
John Guillermin	http://en.wikipedia.org/wiki/John_Guillermin
John Gunther	http://en.wikipedia.org/wiki/John_Gunther
John H. Bryan	http://en.wikipedia.org/wiki/John_H._Bryan
John H. Chafee	http://en.wikipedia.org/wiki/John_H._Chafee
John H. Chafee	http://en.wikipedia.org/wiki/John_H._Chafee
John H. Dalton	http://en.wikipedia.org/wiki/John_H._Dalton
John H. Glenn Jr.	http://en.wikipedia.org/wiki/John_H._Glenn_Jr.
John H. Kinkead	http://en.wikipedia.org/wiki/John_H._Kinkead
John H. Northrop	http://en.wikipedia.org/wiki/John_H._Northrop
John H. Sununu	http://en.wikipedia.org/wiki/John_H._Sununu
John H. Tyson	http://en.wikipedia.org/wiki/John_H._Tyson
John H. van Vleck	http://en.wikipedia.org/wiki/John_H._van_Vleck
John Hall	http://en.wikipedia.org/wiki/John_Hall_(US_politician)
John Hampden	http://en.wikipedia.org/wiki/John_Hampden
John Hancock	http://en.wikipedia.org/wiki/John_Hancock
John Hannah	http://en.wikipedia.org/wiki/John_Hannah_(actor)
John Hannah	http://en.wikipedia.org/wiki/John_Hannah_(American_football)
John Hannah	http://en.wikipedia.org/wiki/John_Hannah_(actor)
John Hanson	http://en.wikipedia.org/wiki/John_Hanson
John Harrison	http://en.wikipedia.org/wiki/John_Harrison
John Hart	http://en.wikipedia.org/wiki/John_Hart
John Hart Ely	http://en.wikipedia.org/wiki/John_Hart_Ely
John Harvard	http://en.wikipedia.org/wiki/John_Harvard_(clergyman)
John Harwood	http://en.wikipedia.org/wiki/John_Harwood
John Hawkes	http://en.wikipedia.org/wiki/John_Hawkes_(actor)
John Hawkes	http://en.wikipedia.org/wiki/John_Hawkes_(novelist)
John Hawkesworth	http://en.wikipedia.org/wiki/John_Hawkesworth_(book_editor)
John Hay	http://en.wikipedia.org/wiki/John_Hay
John Hay Whitney	http://en.wikipedia.org/wiki/John_Hay_Whitney
John Hayes	http://en.wikipedia.org/wiki/John_Henry_Hayes
John Healey	http://en.wikipedia.org/wiki/John_Healey
John Heard	http://en.wikipedia.org/wiki/John_Heard_(actor)
John Heinz	http://en.wikipedia.org/wiki/John_Heinz
John Heinz	http://en.wikipedia.org/wiki/John_Heinz
John Hemming	http://en.wikipedia.org/wiki/John_Hemming_(politician)
John Hench	http://en.wikipedia.org/wiki/John_Hench
John Henry Newman	http://en.wikipedia.org/wiki/John_Henry_Newman
John Hensley	http://en.wikipedia.org/wiki/John_Hensley
John Henson	http://en.wikipedia.org/wiki/John_Henson
John Herschel	http://en.wikipedia.org/wiki/John_Herschel
John Hersey	http://en.wikipedia.org/wiki/John_Hersey
John Hewitt	http://en.wikipedia.org/wiki/John_Hewitt_(poet)
John Heywood	http://en.wikipedia.org/wiki/John_Heywood
John Hiler	http://en.wikipedia.org/wiki/John_Hiler
John Hillerman	http://en.wikipedia.org/wiki/John_Hillerman
John Hinckley	http://en.wikipedia.org/wiki/John_Hinckley
John Hodgman	http://en.wikipedia.org/wiki/John_Hodgman
John Hodiak	http://en.wikipedia.org/wiki/John_Hodiak
John Hoeven	http://en.wikipedia.org/wiki/John_Hoeven
John Hoeven	http://en.wikipedia.org/wiki/John_Hoeven
John Hollander	http://en.wikipedia.org/wiki/John_Hollander
John Holmes	http://en.wikipedia.org/wiki/John_Holmes_(actor)
John Home	http://en.wikipedia.org/wiki/John_Home
John Hooper	http://en.wikipedia.org/wiki/John_Hooper
John Hope Franklin	http://en.wikipedia.org/wiki/John_Hope_Franklin
John Hopkinson	http://en.wikipedia.org/wiki/John_Hopkinson
John Hoppner	http://en.wikipedia.org/wiki/John_Hoppner
John Horrocks	http://en.wikipedia.org/wiki/John_Horrocks_(cotton_manufacturer)
John Hospers	http://en.wikipedia.org/wiki/John_Hospers
John Hostettler	http://en.wikipedia.org/wiki/John_Hostettler
John Houseman	http://en.wikipedia.org/wiki/John_Houseman
John Howard	http://en.wikipedia.org/wiki/John_Howard
John Howard	http://en.wikipedia.org/wiki/John_Howard
John Howard	http://en.wikipedia.org/wiki/John_Howard
John Howard	http://en.wikipedia.org/wiki/John_Howard
John Howard Lawson	http://en.wikipedia.org/wiki/John_Howard_Lawson
John Howe	http://en.wikipedia.org/wiki/John_Howe_(Puritan)
John Howell	http://en.wikipedia.org/wiki/John_Howell_(politician)
John Hughes	http://en.wikipedia.org/wiki/John_Hughes_(filmmaker)
John Hume	http://en.wikipedia.org/wiki/John_Hume
John Hunter	http://en.wikipedia.org/wiki/John_Hunter_(surgeon)
John Hurt	http://en.wikipedia.org/wiki/John_Hurt
John Huston	http://en.wikipedia.org/wiki/John_Huston
John I Tzimisces	http://en.wikipedia.org/wiki/John_I_Tzimisces
John II Comnenus	http://en.wikipedia.org/wiki/John_II_Comnenus
John III Ducas Vatatzes	http://en.wikipedia.org/wiki/John_III_Ducas_Vatatzes
John III Sobieski	http://en.wikipedia.org/wiki/John_III_Sobieski
John Inman	http://en.wikipedia.org/wiki/John_Inman
John Ireland	http://en.wikipedia.org/wiki/John_Ireland_(actor)
John Irving	http://en.wikipedia.org/wiki/John_Irving
John J. Duncan, Sr.	http://en.wikipedia.org/wiki/John_J._Duncan%2C_Sr.
John J. Hamre	http://en.wikipedia.org/wiki/John_J._Hamre
John J. LaFalce	http://en.wikipedia.org/wiki/John_J._LaFalce
John J. McCloy	http://en.wikipedia.org/wiki/John_J._McCloy
John J. O'Connor III	http://en.wikipedia.org/wiki/John_J._O%27Connor_III
John J. Pershing	http://en.wikipedia.org/wiki/John_J._Pershing
John J. Raskob	http://en.wikipedia.org/wiki/John_J._Raskob
John Jacob Astor	http://en.wikipedia.org/wiki/John_Jacob_Astor
John James Audubon	http://en.wikipedia.org/wiki/John_James_Audubon
John Jay	http://en.wikipedia.org/wiki/John_Jay
John Jewel	http://en.wikipedia.org/wiki/John_Jewel
John Joseph Moakley	http://en.wikipedia.org/wiki/John_Joseph_Moakley
John Kander	http://en.wikipedia.org/wiki/John_Kander
John Karlen	http://en.wikipedia.org/wiki/John_Karlen
John Kasich	http://en.wikipedia.org/wiki/John_Kasich
John Keats	http://en.wikipedia.org/wiki/John_Keats
John Kennedy Toole	http://en.wikipedia.org/wiki/John_Kennedy_Toole
John Kenneth Galbraith	http://en.wikipedia.org/wiki/John_Kenneth_Galbraith
John Kerry	http://en.wikipedia.org/wiki/John_Kerry
John Key	http://en.wikipedia.org/wiki/John_Key
John Kitzhaber	http://en.wikipedia.org/wiki/John_Kitzhaber
John Kline	http://en.wikipedia.org/wiki/John_Kline_(politician)
John Kluge	http://en.wikipedia.org/wiki/John_Kluge
John Knowles	http://en.wikipedia.org/wiki/John_Knowles
John Knox	http://en.wikipedia.org/wiki/John_Knox
John Kricfalusi	http://en.wikipedia.org/wiki/John_Kricfalusi
John Kufuor	http://en.wikipedia.org/wiki/John_Kufuor
John L. Burton	http://en.wikipedia.org/wiki/John_L._Burton
John Landis	http://en.wikipedia.org/wiki/John_Landis
John Langdon	http://en.wikipedia.org/wiki/John_Langdon
John Larroquette	http://en.wikipedia.org/wiki/John_Larroquette
John Larson	http://en.wikipedia.org/wiki/John_Larson
John Lasseter	http://en.wikipedia.org/wiki/John_Lasseter
John Latsis	http://en.wikipedia.org/wiki/John_Latsis
John Laurens	http://en.wikipedia.org/wiki/John_Laurens
John Le Carr�	http://en.wikipedia.org/wiki/John_Le_Carr%C3%A9
John Le Mesurier	http://en.wikipedia.org/wiki/John_Le_Mesurier
John Ledyard	http://en.wikipedia.org/wiki/John_Ledyard
John Lee Hooker	http://en.wikipedia.org/wiki/John_Lee_Hooker
John Leech	http://en.wikipedia.org/wiki/John_Leech_(politician)
John Leeson	http://en.wikipedia.org/wiki/John_Leeson
John Legend	http://en.wikipedia.org/wiki/John_Legend
John Leguizamo	http://en.wikipedia.org/wiki/John_Leguizamo
John Lehmann	http://en.wikipedia.org/wiki/John_Lehmann
John Lennon	http://en.wikipedia.org/wiki/John_Lennon
John Lewis	http://en.wikipedia.org/wiki/John_Lewis_(U.S._politician)
John Linder	http://en.wikipedia.org/wiki/John_Linder
John Linnell	http://en.wikipedia.org/wiki/John_Linnell
John Litel	http://en.wikipedia.org/wiki/John_Litel
John Lithgow	http://en.wikipedia.org/wiki/John_Lithgow
John Lloyd Stephens	http://en.wikipedia.org/wiki/John_Lloyd_Stephens
John Locke	http://en.wikipedia.org/wiki/John_Locke
John Lothrop Motley	http://en.wikipedia.org/wiki/John_Lothrop_Motley
John Loudon McAdam	http://en.wikipedia.org/wiki/John_Loudon_McAdam
John Lund	http://en.wikipedia.org/wiki/John_Lund
John Lurie	http://en.wikipedia.org/wiki/John_Lurie
John Lyly	http://en.wikipedia.org/wiki/John_Lyly
John Lynch	http://en.wikipedia.org/wiki/John_Lynch_(New_Hampshire)
John Lynch	http://en.wikipedia.org/wiki/John_Lynch_(New_Hampshire)
John Lynch	http://en.wikipedia.org/wiki/John_Lynch_(actor)
John M. Ford	http://en.wikipedia.org/wiki/John_M._Ford
John M. McConnell	http://en.wikipedia.org/wiki/John_M._McConnell
John M. Murphy	http://en.wikipedia.org/wiki/John_M._Murphy
John M. Spratt, Jr.	http://en.wikipedia.org/wiki/John_M._Spratt%2C_Jr.
John MacArthur	http://en.wikipedia.org/wiki/John_F._MacArthur
John Mack	http://en.wikipedia.org/wiki/John_Edward_Mack
John Madden	http://en.wikipedia.org/wiki/John_Madden_(American_football)
John Mahoney	http://en.wikipedia.org/wiki/John_Mahoney
John Major	http://en.wikipedia.org/wiki/John_Major
John Malkovich	http://en.wikipedia.org/wiki/John_Malkovich
John Mann	http://en.wikipedia.org/wiki/John_Mann_(politician)
John Markoff	http://en.wikipedia.org/wiki/John_Markoff
John Marshall	http://en.wikipedia.org/wiki/John_Marshall
John Marshall Harlan	http://en.wikipedia.org/wiki/John_Marshall_Harlan
John Masefield	http://en.wikipedia.org/wiki/John_Masefield
John Maxwell Coetzee	http://en.wikipedia.org/wiki/John_Maxwell_Coetzee
John Mayall	http://en.wikipedia.org/wiki/John_Mayall
John Mayer	http://en.wikipedia.org/wiki/John_Mayer
John Maynard Keynes	http://en.wikipedia.org/wiki/John_Maynard_Keynes
John Maynard Smith	http://en.wikipedia.org/wiki/John_Maynard_Smith
John McAfee	http://en.wikipedia.org/wiki/John_McAfee
John McAllister Schofield	http://en.wikipedia.org/wiki/John_McAllister_Schofield
John McCain	http://en.wikipedia.org/wiki/John_McCain
John McCarthy	http://en.wikipedia.org/wiki/John_McCarthy_(computer_scientist)
John McCone	http://en.wikipedia.org/wiki/John_McCone
John McDonnell	http://en.wikipedia.org/wiki/John_McDonnell_(politician)
John McDouall Stuart	http://en.wikipedia.org/wiki/John_McDouall_Stuart
John McEnroe	http://en.wikipedia.org/wiki/John_McEnroe
John McEntire	http://en.wikipedia.org/wiki/John_McEntire
John McGahern	http://en.wikipedia.org/wiki/John_McGahern
John McGeoch	http://en.wikipedia.org/wiki/John_McGeoch
John McGraw	http://en.wikipedia.org/wiki/John_McGraw
John McHugh	http://en.wikipedia.org/wiki/John_M._McHugh
John McLaughlin	http://en.wikipedia.org/wiki/John_McLaughlin_(musician)
John McLaughlin	http://en.wikipedia.org/wiki/John_McLaughlin_(host)
John McNaughton	http://en.wikipedia.org/wiki/John_McNaughton
John McPhee	http://en.wikipedia.org/wiki/John_McPhee
John McTiernan	http://en.wikipedia.org/wiki/John_McTiernan
John McVie	http://en.wikipedia.org/wiki/John_McVie
John Melcher	http://en.wikipedia.org/wiki/John_Melcher
John Mica	http://en.wikipedia.org/wiki/John_Mica
John Michell	http://en.wikipedia.org/wiki/John_Michell
John Middleton Clayton	http://en.wikipedia.org/wiki/John_Middleton_Clayton
John Middleton Murry	http://en.wikipedia.org/wiki/John_Middleton_Murry
John Milius	http://en.wikipedia.org/wiki/John_Milius
John Miller	http://en.wikipedia.org/wiki/John_Miller_(Washington)
John Millington Synge	http://en.wikipedia.org/wiki/John_Millington_Synge
John Mills	http://en.wikipedia.org/wiki/John_Mills
John Mills-Cockell	http://en.wikipedia.org/wiki/John_Mills-Cockell
John Milton	http://en.wikipedia.org/wiki/John_Milton
John Mitchell	http://en.wikipedia.org/wiki/John_N._Mitchell
John Mortimer	http://en.wikipedia.org/wiki/John_Mortimer
John Motson	http://en.wikipedia.org/wiki/John_Motson
John Muir	http://en.wikipedia.org/wiki/John_Muir
John N. Dalton	http://en.wikipedia.org/wiki/John_N._Dalton
John Nance Garner	http://en.wikipedia.org/wiki/John_Nance_Garner
John Nash	http://en.wikipedia.org/wiki/John_Forbes_Nash,_Jr.
John Nash	http://en.wikipedia.org/wiki/John_Nash_(architect)
John Neal	http://en.wikipedia.org/wiki/John_Neal
John Negroponte	http://en.wikipedia.org/wiki/John_Negroponte
John Newton	http://en.wikipedia.org/wiki/John_Newton
John Newton	http://en.wikipedia.org/wiki/John_Newton
John Norman	http://en.wikipedia.org/wiki/John_Norman
John Oates	http://en.wikipedia.org/wiki/John_Oates
John Oecolampadius	http://en.wikipedia.org/wiki/John_Oecolampadius
John of Damascus	http://en.wikipedia.org/wiki/John_of_Damascus
John of Gaunt	http://en.wikipedia.org/wiki/John_of_gaunt
John of Salisbury	http://en.wikipedia.org/wiki/John_of_Salisbury
John Ogilby	http://en.wikipedia.org/wiki/John_Ogilby
John O'Hara	http://en.wikipedia.org/wiki/John_O%27Hara
John O'Hurley	http://en.wikipedia.org/wiki/John_O%27Hurley
John Olver	http://en.wikipedia.org/wiki/John_Olver
John Opie	http://en.wikipedia.org/wiki/John_Opie
John Osborne	http://en.wikipedia.org/wiki/John_Osborne
John P. East	http://en.wikipedia.org/wiki/John_P._East
John P. Marquand	http://en.wikipedia.org/wiki/John_P._Marquand
John P. Murtha	http://en.wikipedia.org/wiki/John_Murtha
John Pankow	http://en.wikipedia.org/wiki/John_Pankow
John Parker Hale	http://en.wikipedia.org/wiki/John_Parker_Hale
John Paul Hammerschmidt	http://en.wikipedia.org/wiki/John_Paul_Hammerschmidt
John Paul I	http://en.wikipedia.org/wiki/John_Paul_I
John Paul II	http://en.wikipedia.org/wiki/John_Paul_II
John Paul Jones	http://en.wikipedia.org/wiki/John_Paul_Jones_(musician)
John Paul Jones	http://en.wikipedia.org/wiki/John_Paul_Jones
John Paul Stevens	http://en.wikipedia.org/wiki/John_Paul_Stevens
John Payne	http://en.wikipedia.org/wiki/John_Payne_(actor)
John Peel	http://en.wikipedia.org/wiki/John_peel
John Pendleton Kennedy	http://en.wikipedia.org/wiki/John_Pendleton_Kennedy
John Penrose	http://en.wikipedia.org/wiki/John_Penrose_(politician)
John Perkins	http://en.wikipedia.org/wiki/John_Perkins_(author)
John Perry Barlow	http://en.wikipedia.org/wiki/John_Perry_Barlow
John Peter Altgeld	http://en.wikipedia.org/wiki/John_Peter_Altgeld
John Peterson	http://en.wikipedia.org/wiki/John_E._Peterson
John Petrucci	http://en.wikipedia.org/wiki/John_Petrucci
John Philip Sousa	http://en.wikipedia.org/wiki/John_Philip_Sousa
John Philips	http://en.wikipedia.org/wiki/John_Philips
John Phillip Law	http://en.wikipedia.org/wiki/John_Phillip_Law
John Phillips	http://en.wikipedia.org/wiki/John_Phillips_(musician)
John Philp Thompson	http://en.wikipedia.org/wiki/John_Philp_Thompson,_Sr.
John Playfair	http://en.wikipedia.org/wiki/John_Playfair
John Podesta	http://en.wikipedia.org/wiki/John_Podesta
John Podhoretz	http://en.wikipedia.org/wiki/John_Podhoretz
John Poindexter	http://en.wikipedia.org/wiki/John_Poindexter
John Pope	http://en.wikipedia.org/wiki/John_Pope_(military_officer)
John Popper	http://en.wikipedia.org/wiki/John_Popper
John Power	http://en.wikipedia.org/wiki/John_Power
John Profumo	http://en.wikipedia.org/wiki/John_Profumo
John Pugh	http://en.wikipedia.org/wiki/John_Pugh
John Qualen	http://en.wikipedia.org/wiki/John_Qualen
John Quincy Adams	http://en.wikipedia.org/wiki/John_Quincy_Adams
John R. Block	http://en.wikipedia.org/wiki/John_Rusling_Block
John R. Hicks	http://en.wikipedia.org/wiki/John_Hicks
John R. Kasich	http://en.wikipedia.org/wiki/John_R._Kasich
John R. McKernan, Jr.	http://en.wikipedia.org/wiki/John_R._McKernan,_Jr.
John R. Mott	http://en.wikipedia.org/wiki/John_R._Mott
John R. Steelman	http://en.wikipedia.org/wiki/John_R._Steelman
John Ramsey	http://en.wikipedia.org/wiki/John_Bennett_Ramsey
John Randall	http://en.wikipedia.org/wiki/John_Randall_(UK_politician)
John Randolph	http://en.wikipedia.org/wiki/John_Randolph_(actor)
John Ratzenberger	http://en.wikipedia.org/wiki/John_Ratzenberger
John Rechy	http://en.wikipedia.org/wiki/John_Rechy
John Redwood	http://en.wikipedia.org/wiki/John_Redwood
John Reed	http://en.wikipedia.org/wiki/John_Reed_(journalist)
John Rhys-Davies	http://en.wikipedia.org/wiki/John_Rhys-Davies
John Ritter	http://en.wikipedia.org/wiki/John_Ritter
John Robbins	http://en.wikipedia.org/wiki/John_Robbins_(author)
John Robertson	http://en.wikipedia.org/wiki/John_Robertson_(Glasgow_politician)
John Roebling	http://en.wikipedia.org/wiki/John_Roebling
John Romero	http://en.wikipedia.org/wiki/John_Romero
John Romita, Jr.	http://en.wikipedia.org/wiki/John_Romita,_Jr.
John Romita, Sr.	http://en.wikipedia.org/wiki/John_Romita,_Sr.
John Rowland	http://en.wikipedia.org/wiki/John_G._Rowland
John Ruskin	http://en.wikipedia.org/wiki/John_Ruskin
John Russell	http://en.wikipedia.org/wiki/John_Russell_(actor)
John S. Cooper	http://en.wikipedia.org/wiki/John_S._Cooper
John S. McCain III	http://en.wikipedia.org/wiki/John_McCain
John S. Monagan	http://en.wikipedia.org/wiki/John_S._Monagan
John Salazar	http://en.wikipedia.org/wiki/John_Salazar
John Sarbanes	http://en.wikipedia.org/wiki/John_Sarbanes
John Savage	http://en.wikipedia.org/wiki/John_Savage_(actor)
John Saxon	http://en.wikipedia.org/wiki/John_Saxon_(actor)
John Sayles	http://en.wikipedia.org/wiki/John_Sayles
John Schlesinger	http://en.wikipedia.org/wiki/John_Schlesinger
John Schneider	http://en.wikipedia.org/wiki/John_Schneider_(television_actor)
John Schuck	http://en.wikipedia.org/wiki/John_Schuck
John Scott Haldane	http://en.wikipedia.org/wiki/John_Scott_Haldane
John Sculley	http://en.wikipedia.org/wiki/John_Sculley
John Searle	http://en.wikipedia.org/wiki/John_Searle
John Sebastian	http://en.wikipedia.org/wiki/John_Sebastian
John Selden	http://en.wikipedia.org/wiki/John_Selden
John Shadegg	http://en.wikipedia.org/wiki/John_Shadegg
John Shalikashvili	http://en.wikipedia.org/wiki/John_Shalikashvili
John Shelby Spong	http://en.wikipedia.org/wiki/John_Shelby_Spong
John Sherman	http://en.wikipedia.org/wiki/John_Sherman_(politician)
John Shimkus	http://en.wikipedia.org/wiki/John_Shimkus
John Silber	http://en.wikipedia.org/wiki/John_Silber
John Simon	http://en.wikipedia.org/wiki/John_Simon_(critic)
John Singer Sargent	http://en.wikipedia.org/wiki/John_Singer_Sargent
John Singleton	http://en.wikipedia.org/wiki/John_Singleton
John Singleton Copley	http://en.wikipedia.org/wiki/John_Singleton_Copley
John Skelton	http://en.wikipedia.org/wiki/John_Skelton
John Smith	http://en.wikipedia.org/wiki/John_Smith_(explorer)
John Snow	http://en.wikipedia.org/wiki/John_W._Snow
John Spellar	http://en.wikipedia.org/wiki/John_Spellar
John Spencer	http://en.wikipedia.org/wiki/John_Spencer_(actor)
John Spratt	http://en.wikipedia.org/wiki/John_Spratt
John Stamos	http://en.wikipedia.org/wiki/John_Stamos
John Standing	http://en.wikipedia.org/wiki/John_Standing
John Stanley	http://en.wikipedia.org/wiki/John_Stanley_(politician)
John Steinbeck	http://en.wikipedia.org/wiki/John_steinbeck
John Stevens	http://en.wikipedia.org/wiki/John_Stevens_(drummer)
John Stevenson	http://en.wikipedia.org/wiki/John_Stevenson_(UK_politician)
John Stossel	http://en.wikipedia.org/wiki/John_Stossel
John Stow	http://en.wikipedia.org/wiki/John_Stow
John Stuart Mill	http://en.wikipedia.org/wiki/John_Stuart_Mill
John Stuart, 3rd Earl of Bute	http://en.wikipedia.org/wiki/John_Stuart,_3rd_Earl_of_Bute
John Sturges	http://en.wikipedia.org/wiki/John_Sturges
John Sullivan	http://en.wikipedia.org/wiki/John_Sullivan_(U.S._Rep)
John Sullivan	http://en.wikipedia.org/wiki/John_Sullivan
John Sweeney	http://en.wikipedia.org/wiki/John_E._Sweeney
John T. Chambers	http://en.wikipedia.org/wiki/John_T._Chambers
John T. Dunlop	http://en.wikipedia.org/wiki/John_Thomas_Dunlop
John T. Flynn	http://en.wikipedia.org/wiki/John_T._Flynn
John T. Myers	http://en.wikipedia.org/wiki/John_T._Myers_(Congressman)
John T. Walton	http://en.wikipedia.org/wiki/John_T._Walton
John Tanner	http://en.wikipedia.org/wiki/John_Tanner_(U.S._Representative)
John Tayler	http://en.wikipedia.org/wiki/John_Tayler
John Taylor	http://en.wikipedia.org/wiki/John_Taylor_(bass_guitarist)
John Taylor	http://en.wikipedia.org/wiki/John_Taylor_(poet)
John Terry	http://en.wikipedia.org/wiki/John_Terry
John Tesh	http://en.wikipedia.org/wiki/John_Tesh
John Thaw	http://en.wikipedia.org/wiki/John_Thaw
John the Baptist	http://en.wikipedia.org/wiki/John_the_baptist
John Thompson	http://en.wikipedia.org/wiki/John_Sparrow_David_Thompson
John Thune	http://en.wikipedia.org/wiki/John_Thune
John Thurso	http://en.wikipedia.org/wiki/John_Thurso
John Tierney	http://en.wikipedia.org/wiki/John_F._Tierney
John Toland	http://en.wikipedia.org/wiki/John_Toland_(author)
John Torrey	http://en.wikipedia.org/wiki/John_Torrey
John Tower	http://en.wikipedia.org/wiki/John_Tower
John Travolta	http://en.wikipedia.org/wiki/John_travolta
John Trumbull	http://en.wikipedia.org/wiki/John_Trumbull
John Turner	http://en.wikipedia.org/wiki/John_Turner
John Turturro	http://en.wikipedia.org/wiki/John_Turturro
John Tyler	http://en.wikipedia.org/wiki/John_tyler
John Updike	http://en.wikipedia.org/wiki/John_Updike
John Vanbrugh	http://en.wikipedia.org/wiki/John_Vanbrugh
John Vanderlyn	http://en.wikipedia.org/wiki/John_Vanderlyn
John Varley	http://en.wikipedia.org/wiki/John_Varley_(author)
John Ventimiglia	http://en.wikipedia.org/wiki/John_Ventimiglia
John Vernon	http://en.wikipedia.org/wiki/John_Vernon
John Vessey	http://en.wikipedia.org/wiki/John_Vessey
John von Neumann	http://en.wikipedia.org/wiki/John_von_neumann
John W. Jenrette, Jr.	http://en.wikipedia.org/wiki/John_Jenrette
John W. Seybold	http://en.wikipedia.org/wiki/John_W._Seybold
John W. Thompson	http://en.wikipedia.org/wiki/John_W._Thompson
John W. Troy	http://en.wikipedia.org/wiki/John_Weir_Troy
John W. Warner	http://en.wikipedia.org/wiki/John_Warner
John Waite	http://en.wikipedia.org/wiki/John_Waite
John Walker Lindh	http://en.wikipedia.org/wiki/John_Walker_Lindh
John Wallis	http://en.wikipedia.org/wiki/John_wallis
John Walsh	http://en.wikipedia.org/wiki/John_Walsh
John Walters	http://en.wikipedia.org/wiki/John_P._Walters
John Warner	http://en.wikipedia.org/wiki/John_Warner
John Warnock	http://en.wikipedia.org/wiki/John_Warnock
John Waters	http://en.wikipedia.org/wiki/John_Waters_(filmmaker)
John Watson	http://en.wikipedia.org/wiki/John_B._Watson
John Wayne	http://en.wikipedia.org/wiki/John_wayne
John Wayne Bobbitt	http://en.wikipedia.org/wiki/John_Wayne_Bobbitt 
John Wayne Gacy	http://en.wikipedia.org/wiki/John_Wayne_Gacy
John Webster	http://en.wikipedia.org/wiki/John_Webster
John Wesley	http://en.wikipedia.org/wiki/John_Wesley
John Wesley Powell	http://en.wikipedia.org/wiki/John_Wesley_Powell
John Wesley Shipp	http://en.wikipedia.org/wiki/John_Wesley_Shipp
John Wetton	http://en.wikipedia.org/wiki/John_Wetton
John Whitehead	http://en.wikipedia.org/wiki/John_Whitehead_(singer)
John Whittingdale	http://en.wikipedia.org/wiki/John_Whittingdale
John Wickham	http://en.wikipedia.org/wiki/John_A._Wickham,_Jr.
John Wiese	http://en.wikipedia.org/wiki/John_Wiese
John Wilkes	http://en.wikipedia.org/wiki/John_Wilkes
John Wilkes Booth	http://en.wikipedia.org/wiki/John_wilkes_booth
John Wilkins	http://en.wikipedia.org/wiki/John_Wilkins
John William Dawson	http://en.wikipedia.org/wiki/John_William_Dawson
John William Waterhouse	http://en.wikipedia.org/wiki/John_William_Waterhouse
John Williams	http://en.wikipedia.org/wiki/John_williams
John Wilmot	http://en.wikipedia.org/wiki/John_Wilmot,_2nd_Earl_of_Rochester
John Winthrop	http://en.wikipedia.org/wiki/John_Winthrop
John Winthrop the Younger	http://en.wikipedia.org/wiki/John_Winthrop_the_Younger
John Wise	http://en.wikipedia.org/wiki/John_Wise_(clergyman)
John Wojtowicz	http://en.wikipedia.org/wiki/John_Wojtowicz
John Woo	http://en.wikipedia.org/wiki/John_woo
John Woodcock	http://en.wikipedia.org/wiki/John_Woodcock_(UK_politician)
John Wooden	http://en.wikipedia.org/wiki/John_Wooden
John Woolman	http://en.wikipedia.org/wiki/John_Woolman
John Wozniak	http://en.wikipedia.org/wiki/John_Wozniak
John Wycliffe	http://en.wikipedia.org/wiki/John_wycliffe
John Wyndham	http://en.wikipedia.org/wiki/John_Wyndham
John Yarmuth	http://en.wikipedia.org/wiki/John_Yarmuth
John Yoo	http://en.wikipedia.org/wiki/John_Yoo
John Young	http://en.wikipedia.org/wiki/John_Young_(governor)
John Zachary Young	http://en.wikipedia.org/wiki/John_Zachary_Young
John Zarrella	http://en.wikipedia.org/wiki/John_Zarrella
John Zorn	http://en.wikipedia.org/wiki/John_zorn
Johnathon Schaech	http://en.wikipedia.org/wiki/Johnathan_Schaech
Johnnie Cochran	http://en.wikipedia.org/wiki/Johnnie_Cochran
Johnnie Ray	http://en.wikipedia.org/wiki/Johnnie_Ray
Johnny B.	http://en.wikipedia.org/wiki/John_G._Brennan
Johnny Ball	http://en.wikipedia.org/wiki/Johnny_Ball
Johnny Bench	http://en.wikipedia.org/wiki/Johnny_Bench
Johnny Burnette	http://en.wikipedia.org/wiki/Johnny_Burnette
Johnny Carson	http://en.wikipedia.org/wiki/Johnny_carson
Johnny Cash	http://en.wikipedia.org/wiki/Johnny_cash
Johnny Crawford	http://en.wikipedia.org/wiki/Johnny_Crawford
Johnny Damon	http://en.wikipedia.org/wiki/Johnny_Damon
Johnny Depp	http://en.wikipedia.org/wiki/Johnny_depp
Johnny Galecki	http://en.wikipedia.org/wiki/Johnny_Galecki
Johnny Gill	http://en.wikipedia.org/wiki/Johnny_Gill
Johnny Hallyday	http://en.wikipedia.org/wiki/Johnny_Hallyday
Johnny Hart	http://en.wikipedia.org/wiki/Johnny_Hart
Johnny Isakson	http://en.wikipedia.org/wiki/Johnny_Isakson
Johnny Kelly	http://en.wikipedia.org/wiki/Johnny_Kelly
Johnny Kidd	http://en.wikipedia.org/wiki/Johnny_Kidd_(singer)
Johnny Knoxville	http://en.wikipedia.org/wiki/Johnny_Knoxville
Johnny Mack Brown	http://en.wikipedia.org/wiki/Johnny_Mack_Brown
Johnny Marr	http://en.wikipedia.org/wiki/Johnny_Marr
Johnny Mathis	http://en.wikipedia.org/wiki/Johnny_Mathis
Johnny Mercer	http://en.wikipedia.org/wiki/Johnny_Mercer
Johnny Oates	http://en.wikipedia.org/wiki/Johnny_Oates
Johnny Olson	http://en.wikipedia.org/wiki/Johnny_Olson
Johnny Otis	http://en.wikipedia.org/wiki/Johnny_Otis
Johnny Paycheck	http://en.wikipedia.org/wiki/Johnny_Paycheck
Johnny Ramone	http://en.wikipedia.org/wiki/Johnny_Ramone
Johnny Rebel	http://en.wikipedia.org/wiki/Johnny_Rebel_(singer)
Johnny Rotten	http://en.wikipedia.org/wiki/Johnny_Rotten
Johnny Rutherford	http://en.wikipedia.org/wiki/Johnny_Rutherford
Johnny Rzeznik	http://en.wikipedia.org/wiki/Johnny_Rzeznik
Johnny Thunders	http://en.wikipedia.org/wiki/Johnny_Thunders
Johnny Unitas	http://en.wikipedia.org/wiki/Johnny_Unitas
Johnny Weissmuller	http://en.wikipedia.org/wiki/Johnny_Weissmuller
Johnny Whitworth	http://en.wikipedia.org/wiki/Johnny_Whitworth
Johnny Winter	http://en.wikipedia.org/wiki/Johnny_Winter
Johnson Toribiong	http://en.wikipedia.org/wiki/Johnson_Toribiong
Jolene Blalock	http://en.wikipedia.org/wiki/Jolene_Blalock
Jolin Tsai	http://en.wikipedia.org/wiki/Jolin_Tsai
Jomo Kenyatta	http://en.wikipedia.org/wiki/Jomo_Kenyatta
Jon Anderson	http://en.wikipedia.org/wiki/Jon_Anderson
Jon Avnet	http://en.wikipedia.org/wiki/Jon_Avnet
Jon Bon Jovi	http://en.wikipedia.org/wiki/Jon_Bon_Jovi
Jon Carter	http://en.wikipedia.org/wiki/Jon_Carter
Jon Corzine	http://en.wikipedia.org/wiki/Jon_corzine
Jon Crosby	http://en.wikipedia.org/wiki/Jon_Crosby
Jon Cruddas	http://en.wikipedia.org/wiki/Jon_Cruddas
Jon Cryer	http://en.wikipedia.org/wiki/Jon_Cryer
Jon Favreau	http://en.wikipedia.org/wiki/Jon_Favreau
Jon Fishman	http://en.wikipedia.org/wiki/Jon_Fishman
Jon Hall	http://en.wikipedia.org/wiki/Jon_Hall
Jon Heder	http://en.wikipedia.org/wiki/Jon_Heder
Jon Huntsman, Jr.	http://en.wikipedia.org/wiki/Jon_Huntsman,_Jr.
Jon Johansen	http://en.wikipedia.org/wiki/Jon_Johansen
Jon Krakauer	http://en.wikipedia.org/wiki/Jon_Krakauer
Jon Kyl	http://en.wikipedia.org/wiki/Jon_Kyl
Jon Lovitz	http://en.wikipedia.org/wiki/Jon_Lovitz
Jon Meacham	http://en.wikipedia.org/wiki/Jon_Meacham
Jon Pertwee	http://en.wikipedia.org/wiki/Jon_Pertwee
Jon Polito	http://en.wikipedia.org/wiki/Jon_Polito
Jon Porter	http://en.wikipedia.org/wiki/Jon_Porter
Jon Postel	http://en.wikipedia.org/wiki/Jon_Postel
Jon Provost	http://en.wikipedia.org/wiki/Jon_Provost
Jon Secada	http://en.wikipedia.org/wiki/Jon_Secada
Jon Seda	http://en.wikipedia.org/wiki/Jon_Seda
Jon Stewart	http://en.wikipedia.org/wiki/Jon_stewart
Jon Tester	http://en.wikipedia.org/wiki/Jon_Tester
Jon Trickett	http://en.wikipedia.org/wiki/Jon_Trickett
Jon Turteltaub	http://en.wikipedia.org/wiki/Jon_Turteltaub
Jon Voight	http://en.wikipedia.org/wiki/Jon_voight
Jonah Goldberg	http://en.wikipedia.org/wiki/Jonah_Goldberg
Jonas Salk	http://en.wikipedia.org/wiki/Jonas_Salk
Jonas Savimbi	http://en.wikipedia.org/wiki/Jonas_Savimbi
Jonathan Alter	http://en.wikipedia.org/wiki/Jonathan_Alter
Jonathan Banks	http://en.wikipedia.org/wiki/Jonathan_Banks
Jonathan Brandis	http://en.wikipedia.org/wiki/Jonathan_Brandis
Jonathan Coe	http://en.wikipedia.org/wiki/Jonathan_Coe
Jonathan D. Moreno	http://en.wikipedia.org/wiki/Jonathan_D._Moreno
Jonathan Daniels	http://en.wikipedia.org/wiki/Jonathan_W._Daniels
Jonathan Davis	http://en.wikipedia.org/wiki/Jonathan_Davis
Jonathan Demme	http://en.wikipedia.org/wiki/Jonathan_Demme
Jonathan Djanogly	http://en.wikipedia.org/wiki/Jonathan_Djanogly
Jonathan Edwards	http://en.wikipedia.org/wiki/Jonathan_Edwards_(Welsh_politician)
Jonathan Edwards	http://en.wikipedia.org/wiki/Jonathan_Edwards_(theologian)
Jonathan Evans	http://en.wikipedia.org/wiki/Jonathan_Evans_(politician)
Jonathan Frakes	http://en.wikipedia.org/wiki/Jonathan_Frakes
Jonathan Franzen	http://en.wikipedia.org/wiki/Jonathan_Franzen
Jonathan Frid	http://en.wikipedia.org/wiki/Jonathan_Frid
Jonathan Gilbert	http://en.wikipedia.org/wiki/Jonathan_Gilbert
Jonathan Harris	http://en.wikipedia.org/wiki/Jonathan_Harris
Jonathan J. Bush	http://en.wikipedia.org/wiki/Jonathan_Bush
Jonathan Jackson	http://en.wikipedia.org/wiki/Jonathan_Jackson_(actor)
Jonathan Kaplan	http://en.wikipedia.org/wiki/Jonathan_Kaplan
Jonathan Katz	http://en.wikipedia.org/wiki/Jonathan_Katz
Jonathan King	http://en.wikipedia.org/wiki/Jonathan_King
Jonathan Kozol	http://en.wikipedia.org/wiki/Jonathan_Kozol
Jonathan Lethem	http://en.wikipedia.org/wiki/Jonathan_Lethem
Jonathan Lipnicki	http://en.wikipedia.org/wiki/Jonathan_Lipnicki
Jonathan Lord	http://en.wikipedia.org/wiki/Jonathan_Lord
Jonathan M. Wainwright	http://en.wikipedia.org/wiki/Jonathan_Mayhew_Wainwright_IV
Jonathan Mayhew	http://en.wikipedia.org/wiki/Jonathan_Mayhew
Jonathan Miller	http://en.wikipedia.org/wiki/Jonathan_Miller
Jonathan Pryce	http://en.wikipedia.org/wiki/Jonathan_Pryce
Jonathan Reynolds	http://en.wikipedia.org/wiki/Jonathan_Reynolds
Jonathan Rhys-Meyers	http://en.wikipedia.org/wiki/Jonathan_Rhys_Meyers
Jonathan Richman	http://en.wikipedia.org/wiki/Jonathan_Richman
Jonathan S. Adelstein	http://en.wikipedia.org/wiki/Jonathan_S._Adelstein
Jonathan Segel	http://en.wikipedia.org/wiki/Jonathan_Segel
Jonathan Silverman	http://en.wikipedia.org/wiki/Jonathan_Silverman
Jonathan Swift	http://en.wikipedia.org/wiki/Jonathan_Swift
Jonathan Taylor Thomas	http://en.wikipedia.org/wiki/Jonathan_Taylor_Thomas
Jonathan Turley	http://en.wikipedia.org/wiki/Jonathan_Turley
Jonathan Winters	http://en.wikipedia.org/wiki/Jonathan_Winters
JonBen�t Ramsey	http://en.wikipedia.org/wiki/JonBen�t_Ramsey
Jon-Erik Hexum	http://en.wikipedia.org/wiki/Jon-Erik_Hexum
Jones Very	http://en.wikipedia.org/wiki/Jones_Very
Joni Mitchell	http://en.wikipedia.org/wiki/Joni_Mitchell
Jonny Greenwood	http://en.wikipedia.org/wiki/Jonny_Greenwood
Jonny Lee Miller	http://en.wikipedia.org/wiki/Jonny_Lee_Miller
J�ns Jacob Berzelius	http://en.wikipedia.org/wiki/J�ns_Jacob_Berzelius
Jordan Knight	http://en.wikipedia.org/wiki/Jordan_Knight
Jordana Brewster	http://en.wikipedia.org/wiki/Jordana_Brewster
J�rg Haider	http://en.wikipedia.org/wiki/J�rg_Haider
Jorge Amado	http://en.wikipedia.org/wiki/Jorge_Amado
Jorge Garcia	http://en.wikipedia.org/wiki/Jorge_Garcia
Jorge Luis Borges	http://en.wikipedia.org/wiki/Jorge_Luis_Borges
Jorge Posada	http://en.wikipedia.org/wiki/Jorge_Posada
Jorge Sampaio	http://en.wikipedia.org/wiki/Jorge_Sampaio 
Jorie Graham	http://en.wikipedia.org/wiki/Jorie_Graham
Joris-Karl Huysmans	http://en.wikipedia.org/wiki/Joris-Karl_Huysmans
Jorja Fox	http://en.wikipedia.org/wiki/Jorja_Fox
Joscelyn Godwin	http://en.wikipedia.org/wiki/Joscelyn_Godwin
Joschka Fischer	http://en.wikipedia.org/wiki/Joschka_Fischer
Jos� Agostinho de Macedo	http://en.wikipedia.org/wiki/Jos�_Agostinho_de_Macedo
Jos� Antonio P�ez	http://en.wikipedia.org/wiki/Jos�_Antonio_P�ez
Jose Canseco	http://en.wikipedia.org/wiki/Jose_Canseco
Jos� Carreras	http://en.wikipedia.org/wiki/Jos�_Carreras
Jos� Clemente Orozco	http://en.wikipedia.org/wiki/Jos�_Clemente_Orozco
Jos� de Ribera	http://en.wikipedia.org/wiki/Jusepe_de_Ribera
Jose de San Martin	http://en.wikipedia.org/wiki/Jos�_de_San_Mart�n
Jos� Eber	http://en.wikipedia.org/wiki/Jos�_Eber
Jos� Echegaray	http://en.wikipedia.org/wiki/Jos�_Echegaray
Jos� Eduardo dos Santos	http://en.wikipedia.org/wiki/Jos�_Eduardo_dos_Santos
Jos� Feliciano	http://en.wikipedia.org/wiki/Jos�_Feliciano
Jose Ferrer	http://en.wikipedia.org/wiki/Jos�_Ferrer
Jos� Guadalupe Posada	http://en.wikipedia.org/wiki/Jos�_Guadalupe_Posada
Jos� Luis Rodr�guez Zapatero	http://en.wikipedia.org/wiki/Jos�_Luis_Rodr�guez_Zapatero
Jos� Manuel Barroso	http://en.wikipedia.org/wiki/Dur%C3%A3o_Barroso
Jose Maria Aznar	http://en.wikipedia.org/wiki/Jos�_Mar�a_Aznar
Jos� Mar�a de Heredia	http://en.wikipedia.org/wiki/Jos�-Maria_de_Heredia
Jos� Mar�a de Pereda	http://en.wikipedia.org/wiki/Jos�_Mar�a_de_Pereda
Jose Maria Morelos	http://en.wikipedia.org/wiki/Jos�_Mar�a_Morelos
Jos� Maria Neves	http://en.wikipedia.org/wiki/Jos�_Maria_Neves 
Jos� Mart�nez Ruiz	http://en.wikipedia.org/wiki/Jos�_Mart�nez_Ruiz
Jose Mourinho	http://en.wikipedia.org/wiki/Jos�_Mourinho
Jos� Mujica	http://en.wikipedia.org/wiki/Jos�_Mujica
Jos� Napole�n Duarte	http://en.wikipedia.org/wiki/Jos�_Napole�n_Duarte
Jos� P. Laurel	http://en.wikipedia.org/wiki/Jos�_P._Laurel
Jose Padilla	http://en.wikipedia.org/wiki/Jos�_Padilla_(prisoner)
Jos� Ramos Horta	http://en.wikipedia.org/wiki/Jos�_Ramos-Horta
Jos� Saramago	http://en.wikipedia.org/wiki/Jos�_Saramago
Jos� Serrano	http://en.wikipedia.org/wiki/Jos�_Serrano
Jos� S�crates	http://en.wikipedia.org/wiki/Jos�_S�crates
Josef Albers	http://en.wikipedia.org/wiki/Josef_Albers
Josef Hoffmann	http://en.wikipedia.org/wiki/Josef_Hoffmann
Josef von Sternberg	http://en.wikipedia.org/wiki/Josef_von_Sternberg
Joseph Addison	http://en.wikipedia.org/wiki/Joseph_Addison
Joseph Alioto	http://en.wikipedia.org/wiki/Joseph_Alioto
Joseph Aloysius Hansom	http://en.wikipedia.org/wiki/Joseph_Aloysius_Hansom
Joseph Alsop	http://en.wikipedia.org/wiki/Joseph_Alsop
Joseph Banks Rhine	http://en.wikipedia.org/wiki/Joseph_Banks_Rhine
Joseph Barbera	http://en.wikipedia.org/wiki/Joseph_Barbera
Joseph Beuys	http://en.wikipedia.org/wiki/Joseph_Beuys
Joseph Biden	http://en.wikipedia.org/wiki/Joseph_Biden
Joseph Bologna	http://en.wikipedia.org/wiki/Joseph_Bologna
Joseph Bramah	http://en.wikipedia.org/wiki/Joseph_Bramah
Joseph Brant	http://en.wikipedia.org/wiki/Joseph_Brant
Joseph Brodsky	http://en.wikipedia.org/wiki/Joseph_Brodsky
Joseph C. Yates	http://en.wikipedia.org/wiki/Joseph_C._Yates
Joseph Califano	http://en.wikipedia.org/wiki/Joseph_Califano
Joseph Campanella	http://en.wikipedia.org/wiki/Joseph_Campanella
Joseph Campbell	http://en.wikipedia.org/wiki/Joseph_Campbell
Joseph Cao	http://en.wikipedia.org/wiki/Joseph_Cao
Joseph Chamberlain	http://en.wikipedia.org/wiki/Joseph_Chamberlain
Joseph Conrad	http://en.wikipedia.org/wiki/Joseph_Conrad
Joseph Coors, Sr.	http://en.wikipedia.org/wiki/Joseph_Coors
Joseph Cornell	http://en.wikipedia.org/wiki/Joseph_Cornell
Joseph Cotten	http://en.wikipedia.org/wiki/Joseph_Cotten
Joseph Crowley	http://en.wikipedia.org/wiki/Joseph_Crowley
Joseph D. Early	http://en.wikipedia.org/wiki/Joseph_D._Early
Joseph Dalton Hooker	http://en.wikipedia.org/wiki/Joseph_Dalton_Hooker
Joseph E. Schmitz	http://en.wikipedia.org/wiki/Joseph_E._Schmitz
Joseph Eggleston Johnston	http://en.wikipedia.org/wiki/Joseph_Eggleston_Johnston
Joseph Ejercito Estrada	http://en.wikipedia.org/wiki/Joseph_Ejercito_Estrada
Joseph F. Cullman III	http://en.wikipedia.org/wiki/Joseph_Cullman
Joseph Fiennes	http://en.wikipedia.org/wiki/Joseph_Fiennes
Joseph Glanvill	http://en.wikipedia.org/wiki/Joseph_Glanvill
Joseph Goebbels	http://en.wikipedia.org/wiki/Joseph_Goebbels
Joseph Gordon-Levitt	http://en.wikipedia.org/wiki/Joseph_Gordon-Levitt
Joseph Grew	http://en.wikipedia.org/wiki/Joseph_Grew
Joseph Grimaldi	http://en.wikipedia.org/wiki/Joseph_Grimaldi
Joseph Gurney Cannon	http://en.wikipedia.org/wiki/Joseph_Gurney_Cannon
Joseph H. Himes	http://en.wikipedia.org/wiki/Joseph_H._Himes
Joseph H. Short	http://en.wikipedia.org/wiki/Joseph_H._Short
Joseph H. Taylor, Jr.	http://en.wikipedia.org/wiki/Joseph_H._Taylor
Joseph Hahn	http://en.wikipedia.org/wiki/Joseph_Hahn
Joseph Hall	http://en.wikipedia.org/wiki/Joseph_Hall_(bishop)
Joseph Hansen	http://en.wikipedia.org/wiki/Joseph_Hansen_(writer)
Joseph Haydn	http://en.wikipedia.org/wiki/Joseph_Haydn
Joseph Heller	http://en.wikipedia.org/wiki/Joseph_Heller
Joseph Henry	http://en.wikipedia.org/wiki/Joseph_Henry
Joseph Henry Shorthouse	http://en.wikipedia.org/wiki/Joseph_Henry_Shorthouse
Joseph Hergesheimer	http://en.wikipedia.org/wiki/Joseph_Hergesheimer
Joseph Hoeffel	http://en.wikipedia.org/wiki/Joseph_Hoeffel
Joseph Hooker	http://en.wikipedia.org/wiki/Joseph_Hooker
Joseph Howe	http://en.wikipedia.org/wiki/Joseph_Howe
Joseph I	http://en.wikipedia.org/wiki/Joseph_I,_Holy_Roman_Emperor
Joseph II	http://en.wikipedia.org/wiki/Joseph_II,_Holy_Roman_Emperor
Joseph J. DioGuardi	http://en.wikipedia.org/wiki/Joseph_J._DioGuardi
Joseph Jarman	http://en.wikipedia.org/wiki/Joseph_Jarman
Joseph Joachim	http://en.wikipedia.org/wiki/Joseph_Joachim
Joseph Kabila	http://en.wikipedia.org/wiki/Joseph_Kabila
Joseph Kabui	http://en.wikipedia.org/wiki/Joseph_Kabui
Joseph Kernan	http://en.wikipedia.org/wiki/Joseph_Kernan
Joseph Kirkland	http://en.wikipedia.org/wiki/Joseph_Kirkland
Joseph Knollenberg	http://en.wikipedia.org/wiki/Joseph_Knollenberg
Joseph Konopka	http://en.wikipedia.org/wiki/Joseph_Konopka
Joseph Kony	http://en.wikipedia.org/wiki/Joseph_Kony
Joseph L. Mankiewicz	http://en.wikipedia.org/wiki/Joseph_L._Mankiewicz
Joseph Lieberman	http://en.wikipedia.org/wiki/Joseph_Lieberman
Joseph Lister	http://en.wikipedia.org/wiki/Joseph_Lister,_1st_Baron_Lister
Joseph Losey	http://en.wikipedia.org/wiki/Joseph_Losey
Joseph Lowery	http://en.wikipedia.org/wiki/Joseph_Lowery
Joseph M. Gaydos	http://en.wikipedia.org/wiki/Joseph_M._Gaydos
Joseph M. McDade	http://en.wikipedia.org/wiki/Joseph_M._McDade
Joseph M. Tucci	http://en.wikipedia.org/wiki/Joseph_M._Tucci
Joseph McCarthy	http://en.wikipedia.org/wiki/Joseph_McCarthy
Joseph McElroy	http://en.wikipedia.org/wiki/Joseph_McElroy
Joseph Merrick	http://en.wikipedia.org/wiki/Joseph_Merrick
Joseph Mitchell	http://en.wikipedia.org/wiki/Joseph_Mitchell
Joseph Nacchio	http://en.wikipedia.org/wiki/Joseph_Nacchio
Joseph of Arimathea	http://en.wikipedia.org/wiki/Joseph_of_Arimathea
Joseph P. Addabbo	http://en.wikipedia.org/wiki/Joseph_P._Addabbo
Joseph P. Kennedy	http://en.wikipedia.org/wiki/Joseph_P._Kennedy,_Sr.
Joseph Papp	http://en.wikipedia.org/wiki/Joseph_Papp
Joseph Priestley	http://en.wikipedia.org/wiki/Joseph_Priestley
Joseph Pulitzer	http://en.wikipedia.org/wiki/Joseph_Pulitzer
Joseph R. Biden, Jr.	http://en.wikipedia.org/wiki/Joseph_R._Biden,_Jr.
Joseph R. Pitts	http://en.wikipedia.org/wiki/Joseph_Pitts
Joseph Rotblat	http://en.wikipedia.org/wiki/Joseph_Rotblat
Joseph Sargent	http://en.wikipedia.org/wiki/Joseph_Sargent
Joseph Schildkraut	http://en.wikipedia.org/wiki/Joseph_Schildkraut
Joseph Sill Clark	http://en.wikipedia.org/wiki/Joseph_Sill_Clark
Joseph Smith	http://en.wikipedia.org/wiki/Joseph_Smith,_Jr.
Joseph Stiglitz	http://en.wikipedia.org/wiki/Joseph_Stiglitz
Joseph Stilwell	http://en.wikipedia.org/wiki/Joseph_Stillwell
Joseph Story	http://en.wikipedia.org/wiki/Joseph_Story
Joseph Sturge	http://en.wikipedia.org/wiki/Joseph_Sturge
Joseph Urusemal	http://en.wikipedia.org/wiki/Joseph_Urusemal
Joseph Wambaugh	http://en.wikipedia.org/wiki/Joseph_Wambaugh
Joseph Warren	http://en.wikipedia.org/wiki/Joseph_Warren
Joseph Wilson	http://en.wikipedia.org/wiki/Joseph_C._Wilson
Joseph Wirth	http://en.wikipedia.org/wiki/Joseph_Wirth
Joseph Wood Krutch	http://en.wikipedia.org/wiki/Joseph_Wood_Krutch
Joseph Zito	http://en.wikipedia.org/wiki/Joseph_Zito
Josephine Baker	http://en.wikipedia.org/wiki/Josephine_Baker
Josephine Hart	http://en.wikipedia.org/wiki/Josephine_Hart
Josephine Herbst	http://en.wikipedia.org/wiki/Josephine_Herbst
Josephine Hull	http://en.wikipedia.org/wiki/Josephine_Hull
Josephine Humphreys	http://en.wikipedia.org/wiki/Josephine_Humphreys
Josephine Tey	http://en.wikipedia.org/wiki/Josephine_Tey
Joseph-Louis Gay-Lussac	http://en.wikipedia.org/wiki/Joseph_Louis_Gay-Lussac
Joseph-Louis Lagrange	http://en.wikipedia.org/wiki/Joseph_Louis_Lagrange
Joseph-Marie Jacquard	http://en.wikipedia.org/wiki/Joseph_Marie_Jacquard
Joseph-Nicolas Delisle	http://en.wikipedia.org/wiki/Joseph-Nicolas_Delisle
Josh Billings	http://en.wikipedia.org/wiki/Josh_Billings
Josh Bolten	http://en.wikipedia.org/wiki/Josh_Bolten
Josh Brolin	http://en.wikipedia.org/wiki/Josh_Brolin
Josh Charles	http://en.wikipedia.org/wiki/Josh_Charles
Josh Duhamel	http://en.wikipedia.org/wiki/Josh_Duhamel
Josh Freese	http://en.wikipedia.org/wiki/Josh_Freese
Josh Gibson	http://en.wikipedia.org/wiki/Josh_Gibson
Josh Groban	http://en.wikipedia.org/wiki/Josh_Groban
Josh Hartnett	http://en.wikipedia.org/wiki/Josh_Hartnett
Josh Holloway	http://en.wikipedia.org/wiki/Josh_Holloway
Josh Homme	http://en.wikipedia.org/wiki/Josh_Homme
Josh Lucas	http://en.wikipedia.org/wiki/Josh_Lucas
Josh McDowell	http://en.wikipedia.org/wiki/Josh_McDowell
Josh Peck	http://en.wikipedia.org/wiki/Josh_Peck
Josh Schwartz	http://en.wikipedia.org/wiki/Josh_Schwartz
Josh Silver	http://en.wikipedia.org/wiki/Josh_Silver
Joshua Jackson	http://en.wikipedia.org/wiki/Joshua_Jackson
Joshua Leonard	http://en.wikipedia.org/wiki/Joshua_Leonard
Joshua Micah Marshall	http://en.wikipedia.org/wiki/Joshua_Micah_Marshall
Joshua Reynolds	http://en.wikipedia.org/wiki/Joshua_Reynolds
Joshua Sylvester	http://en.wikipedia.org/wiki/Joshua_Sylvester
Josiah Quincy	http://en.wikipedia.org/wiki/Josiah_Quincy_III
Josiah Wedgwood	http://en.wikipedia.org/wiki/Josiah_Wedgwood
Josias Simmler	http://en.wikipedia.org/wiki/Josias_Simmler
Josip Broz Tito	http://en.wikipedia.org/wiki/Josip_Broz_Tito
Josquin Des Prez	http://en.wikipedia.org/wiki/Josquin_des_Prez
Joss Stone	http://en.wikipedia.org/wiki/Joss_Stone
Joss Whedon	http://en.wikipedia.org/wiki/Joss_Whedon
Jost Amman	http://en.wikipedia.org/wiki/Jost_Amman
Jouett Shouse	http://en.wikipedia.org/wiki/Jouett_Shouse
Joy Behar	http://en.wikipedia.org/wiki/Joy_Behar
Joy Bryant	http://en.wikipedia.org/wiki/Joy_Bryant
Joyce Brothers	http://en.wikipedia.org/wiki/Joyce_Brothers
Joyce Carol Oates	http://en.wikipedia.org/wiki/Joyce_Carol_Oates
Joyce Cary	http://en.wikipedia.org/wiki/Joyce_Cary
Joyce DeWitt	http://en.wikipedia.org/wiki/Joyce_dewitt
Joyce Kilmer	http://en.wikipedia.org/wiki/Joyce_Kilmer
Joyce Meyer	http://en.wikipedia.org/wiki/Joyce_Meyer
Joyce Randolph	http://en.wikipedia.org/wiki/Joyce_Randolph
Joyce Van Patten	http://en.wikipedia.org/wiki/Joyce_Van_Patten
Joycelyn Elders	http://en.wikipedia.org/wiki/Joycelyn_Elders
Jozef Isra�ls	http://en.wikipedia.org/wiki/Jozef_Isra�ls
Jozef Lenart	http://en.wikipedia.org/wiki/Jozef_Len�rt
Juan Antonio Samaranch	http://en.wikipedia.org/wiki/Juan_Antonio_Samaranch
Juan Babauta	http://en.wikipedia.org/wiki/Juan_Babauta
Juan Carlos	http://en.wikipedia.org/wiki/Juan_Carlos_I_of_Spain
Juan Cole	http://en.wikipedia.org/wiki/Juan_Cole
Juan Corona	http://en.wikipedia.org/wiki/Juan_Corona
Juan de Pareja	http://en.wikipedia.org/wiki/Juan_de_Pareja
Juan del Encina	http://en.wikipedia.org/wiki/Juan_del_Encina
Juan Escoiquiz	http://en.wikipedia.org/wiki/Juan_Escoiquiz
Juan Gris	http://en.wikipedia.org/wiki/Juan_Gris
Juan Jos� Ibarretxe Markuartu	http://en.wikipedia.org/wiki/Juan_Jos�_Ibarretxe
Juan Marichal	http://en.wikipedia.org/wiki/Juan_Marichal
Juan Peron	http://en.wikipedia.org/wiki/Juan_Per�n
Juan Ponce de Le�n	http://en.wikipedia.org/wiki/Juan_Ponce_de_Le�n
Juan Ram�n Jim�nez	http://en.wikipedia.org/wiki/Juan_Ram�n_Jim�nez
Juan Trippe	http://en.wikipedia.org/wiki/Juan_Trippe
Juan Williams	http://en.wikipedia.org/wiki/Juan_Williams
Juana de Asbaje	http://en.wikipedia.org/wiki/Juana_de_Asbaje
Juanita M. Kreps	http://en.wikipedia.org/wiki/Juanita_M._Kreps
Juanita Millender-McDonald	http://en.wikipedia.org/wiki/Juanita_Millender-McDonald
Juanita Moore	http://en.wikipedia.org/wiki/Juanita_Moore
Judah ben Samuel Halevi	http://en.wikipedia.org/wiki/Judah_Halevi
Judas Iscariot	http://en.wikipedia.org/wiki/Judas_Iscariot
Judd Apatow	http://en.wikipedia.org/wiki/Judd_Apatow
Judd Gregg	http://en.wikipedia.org/wiki/Judd_Gregg
Judd Hirsch	http://en.wikipedia.org/wiki/Judd_Hirsch
Judd Nelson	http://en.wikipedia.org/wiki/Judd_Nelson
Jude Law	http://en.wikipedia.org/wiki/Jude_Law
Jude Wanniski	http://en.wikipedia.org/wiki/Jude_Wanniski
Judge Joe Brown	http://en.wikipedia.org/wiki/Joe_Brown_(judge)
Judge Judy	http://en.wikipedia.org/wiki/Judith_Sheindlin
Judge Larry Joe	http://en.wikipedia.org/wiki/Larry_Joe_Doherty
Judge Reinhold	http://en.wikipedia.org/wiki/Judge_Reinhold
Judge Wapner	http://en.wikipedia.org/wiki/Joseph_Wapner
Judi Dench	http://en.wikipedia.org/wiki/Judi_Dench
Judith Butler	http://en.wikipedia.org/wiki/Judith_Butler
Judith Ivey	http://en.wikipedia.org/wiki/Judith_Ivey
Judith Jamison	http://en.wikipedia.org/wiki/Judith_Jamison
Judith Krantz	http://en.wikipedia.org/wiki/Judith_Krantz
Judith Leyster	http://en.wikipedia.org/wiki/Judith_Leyster
Judith Light	http://en.wikipedia.org/wiki/Judith_Light
Judith Martin	http://en.wikipedia.org/wiki/Judith_Martin
Judith Miller	http://en.wikipedia.org/wiki/Judith_Miller_(journalist)
Judith O'Dea	http://en.wikipedia.org/wiki/Judith_O'Dea
Judith Reisman	http://en.wikipedia.org/wiki/Judith_Reisman
Judith Wright	http://en.wikipedia.org/wiki/Judith_Wright
Judy Biggert	http://en.wikipedia.org/wiki/Judy_Biggert
Judy Blume	http://en.wikipedia.org/wiki/Judy_Blume
Judy Carne	http://en.wikipedia.org/wiki/Judy_Carne
Judy Chicago	http://en.wikipedia.org/wiki/Judy_Chicago
Judy Chu	http://en.wikipedia.org/wiki/Judy_Chu
Judy Collins	http://en.wikipedia.org/wiki/Judy_Collins
Judy Davis	http://en.wikipedia.org/wiki/Judy_Davis
Judy Garland	http://en.wikipedia.org/wiki/Judy_Garland
Judy Greer	http://en.wikipedia.org/wiki/Judy_Greer
Judy Holliday	http://en.wikipedia.org/wiki/Judy_Holliday
Judy Martz	http://en.wikipedia.org/wiki/Judy_Martz
Judy Norton-Taylor	http://en.wikipedia.org/wiki/Judy_Norton_Taylor
Judy Tyler	http://en.wikipedia.org/wiki/Judy_Tyler
Judy Woodruff	http://en.wikipedia.org/wiki/Judy_Woodruff
Juelz Santana	http://en.wikipedia.org/wiki/Juelz_Santana
Juhan Parts	http://en.wikipedia.org/wiki/Juhan_Parts
Juice Newton	http://en.wikipedia.org/wiki/Juice_Newton
Jules Dassin	http://en.wikipedia.org/wiki/Jules_Dassin
Jules Dupr�	http://en.wikipedia.org/wiki/Jules_Dupr�
Jules Feiffer	http://en.wikipedia.org/wiki/Jules_Feiffer
Jules Gr�vy	http://en.wikipedia.org/wiki/Jules_Gr�vy
Jules Massenet	http://en.wikipedia.org/wiki/Jules_Massenet
Jules Mazarin	http://en.wikipedia.org/wiki/Jules_Mazarin
Jules Michelet	http://en.wikipedia.org/wiki/Jules_Michelet
Jules Shear	http://en.wikipedia.org/wiki/Jules_Shear
Jules Stein	http://en.wikipedia.org/wiki/Jules_Stein
Jules Verne	http://en.wikipedia.org/wiki/Jules_Verne
Julia Barr	http://en.wikipedia.org/wiki/Julia_Barr
Julia Carson	http://en.wikipedia.org/wiki/Julia_Carson
Julia Child	http://en.wikipedia.org/wiki/Julia_Child
Julia Duffy	http://en.wikipedia.org/wiki/Julia_Duffy
Julia Louis-Dreyfus	http://en.wikipedia.org/wiki/Julia_Louis-Dreyfus
Julia Migenes	http://en.wikipedia.org/wiki/Julia_Migenes
Julia Morgan	http://en.wikipedia.org/wiki/Julia_Morgan
Julia Ormond	http://en.wikipedia.org/wiki/Julia_Ormond
Julia Roberts	http://en.wikipedia.org/wiki/Julia_Roberts
Julia Stiles	http://en.wikipedia.org/wiki/Julia_Stiles
Julia Sweeney	http://en.wikipedia.org/wiki/Julia_Sweeney
Julia Volkova	http://en.wikipedia.org/wiki/Yulia_Volkova
Julia Ward Howe	http://en.wikipedia.org/wiki/Julia_Ward_Howe
Julian Amyes	http://en.wikipedia.org/wiki/Julian_Charles_Becket_Amyes
Julian Barnes	http://en.wikipedia.org/wiki/Julian_Barnes
Julian Barratt	http://en.wikipedia.org/wiki/Julian_Barratt
Julian Beck	http://en.wikipedia.org/wiki/Julian_Beck
Julian Bond	http://en.wikipedia.org/wiki/Julian_Bond
Julian Brazier	http://en.wikipedia.org/wiki/Julian_Brazier
Julian C. Dixon	http://en.wikipedia.org/wiki/Julian_C._Dixon
Julian Casablancas	http://en.wikipedia.org/wiki/Julian_Casablancas
Julian Cope	http://en.wikipedia.org/wiki/Julian_Cope
Julian Glover	http://en.wikipedia.org/wiki/Julian_Glover
Julian Grenfell	http://en.wikipedia.org/wiki/Julian_Grenfell
Julian Huppert	http://en.wikipedia.org/wiki/Julian_Huppert
Julian Huxley	http://en.wikipedia.org/wiki/Julian_Huxley
Julian Lennon	http://en.wikipedia.org/wiki/Julian_Lennon
Julian Lewis	http://en.wikipedia.org/wiki/Julian_Lewis
Julian May	http://en.wikipedia.org/wiki/Julian_May
Julian McMahon	http://en.wikipedia.org/wiki/Julian_McMahon
Julian Sands	http://en.wikipedia.org/wiki/Julian_Sands
Julian Schwinger	http://en.wikipedia.org/wiki/Julian_Schwinger
Julian Smith	http://en.wikipedia.org/wiki/Julian_Smith_(politician)
Julian Sturdy	http://en.wikipedia.org/wiki/Julian_Sturdy
Julian the Apostate	http://en.wikipedia.org/wiki/Julian_the_Apostate
Juliana Hatfield	http://en.wikipedia.org/wiki/Juliana_Hatfield
Julianna Margulies	http://en.wikipedia.org/wiki/Julianna_Margulies
Julianne Malveaux	http://en.wikipedia.org/wiki/Julianne_Malveaux
Julianne Moore	http://en.wikipedia.org/wiki/Julianne_Moore
Julianne Nicholson	http://en.wikipedia.org/wiki/Julianne_Nicholson
Julianne Phillips	http://en.wikipedia.org/wiki/Julianne_Phillips
Julie Adams	http://en.wikipedia.org/wiki/Julie_Adams
Julie Andrews	http://en.wikipedia.org/wiki/Julie_Andrews
Julie Bell	http://en.wikipedia.org/wiki/Julie_Bell
Julie Benz	http://en.wikipedia.org/wiki/Julie_Benz
Julie Bishop	http://en.wikipedia.org/wiki/Julie_Bishop_(actress)
Julie Bowen	http://en.wikipedia.org/wiki/Julie_Bowen
Julie Brown	http://en.wikipedia.org/wiki/Julie_Brown
Julie Burchill	http://en.wikipedia.org/wiki/Julie_Burchill
Julie Cafritz	http://en.wikipedia.org/wiki/Julie_Cafritz
Julie Chen	http://en.wikipedia.org/wiki/Julie_Chen
Julie Christie	http://en.wikipedia.org/wiki/Julie_Christie
Julie Delpy	http://en.wikipedia.org/wiki/Julie_Delpy
Julie Doucet	http://en.wikipedia.org/wiki/Julie_Doucet
Julie Elliott	http://en.wikipedia.org/wiki/Julie_Elliott
Julie Hagerty	http://en.wikipedia.org/wiki/Julie_Hagerty
Julie Harris	http://en.wikipedia.org/wiki/Julie_Harris
Julie Hilling	http://en.wikipedia.org/wiki/Julie_Hilling
Julie Kavner	http://en.wikipedia.org/wiki/Julie_Kavner
Julie London	http://en.wikipedia.org/wiki/Julie_London
Julie Newmar	http://en.wikipedia.org/wiki/Julie_Newmar
Julie Nixon Eisenhower	http://en.wikipedia.org/wiki/Julie_Nixon_Eisenhower
Julie Taymor	http://en.wikipedia.org/wiki/Julie_Taymor
Julie Walters	http://en.wikipedia.org/wiki/Julie_Walters
Juliet Mills	http://en.wikipedia.org/wiki/Juliet_Mills
Juliet Prowse	http://en.wikipedia.org/wiki/Juliet_Prowse
Juliet Stevenson	http://en.wikipedia.org/wiki/Juliet_Stevenson
Juliette Binoche	http://en.wikipedia.org/wiki/Juliette_Binoche
Juliette Lewis	http://en.wikipedia.org/wiki/Juliette_Lewis
Julio Cort�zar	http://en.wikipedia.org/wiki/Julio_Cort�zar
Julio Iglesias	http://en.wikipedia.org/wiki/Julio_Iglesias
Julius Axelrod	http://en.wikipedia.org/wiki/Julius_Axelrod
Julius Caesar	http://en.wikipedia.org/wiki/Julius_Caesar
Julius Erving	http://en.wikipedia.org/wiki/Julius_Erving
Julius Nepos	http://en.wikipedia.org/wiki/Julius_Nepos
Julius Robert Mayer	http://en.wikipedia.org/wiki/Julius_Robert_von_Mayer
Julius Rosenberg	http://en.wikipedia.org/wiki/Julius_Rosenberg
Julius Schwartz	http://en.wikipedia.org/wiki/Julius_Schwartz
Julius Streicher	http://en.wikipedia.org/wiki/Julius_Streicher
June Allyson	http://en.wikipedia.org/wiki/June_Allyson
June Carter Cash	http://en.wikipedia.org/wiki/June_Carter_Cash
June Christy	http://en.wikipedia.org/wiki/June_Christy
June Duprez	http://en.wikipedia.org/wiki/June_Duprez
June Foray	http://en.wikipedia.org/wiki/June_Foray
June Haver	http://en.wikipedia.org/wiki/June_Haver
June Havoc	http://en.wikipedia.org/wiki/June_Havoc
June Jordan	http://en.wikipedia.org/wiki/June_Jordan
June Lockhart	http://en.wikipedia.org/wiki/June_Lockhart
June Pointer	http://en.wikipedia.org/wiki/June_Pointer
June Taylor	http://en.wikipedia.org/wiki/June_Taylor
Junichiro Koizumi	http://en.wikipedia.org/wiki/Junichiro_Koizumi
Junior Parker	http://en.wikipedia.org/wiki/Junior_Parker
Junior Walker	http://en.wikipedia.org/wiki/Junior_Walker
Jurelang Zedkaia	http://en.wikipedia.org/wiki/Jurelang_Zedkaia
J�rgen Bartsch	http://en.wikipedia.org/wiki/J�rgen_Bartsch
J�rgen Habermas	http://en.wikipedia.org/wiki/J�rgen_Habermas
Jurgen Klinsmann	http://en.wikipedia.org/wiki/J�rgen_Klinsmann
J�rgen Prochnow	http://en.wikipedia.org/wiki/J�rgen_Prochnow
Jus Addiss	http://en.wikipedia.org/wiki/Jus_Addiss
Justin Berfield	http://en.wikipedia.org/wiki/Justin_Berfield
Justin Bieber	http://en.wikipedia.org/wiki/Justin_Bieber
Justin Chambers	http://en.wikipedia.org/wiki/Justin_Chambers
Justin Chatwin	http://en.wikipedia.org/wiki/Justin_Chatwin
Justin Guarini	http://en.wikipedia.org/wiki/Justin_Guarini
Justin Hawkins	http://en.wikipedia.org/wiki/Justin_Hawkins
Justin Hayward	http://en.wikipedia.org/wiki/Justin_Hayward
Justin Kaplan	http://en.wikipedia.org/wiki/Justin_Kaplan
Justin Kirk	http://en.wikipedia.org/wiki/Justin_Kirk
Justin Lin	http://en.wikipedia.org/wiki/Justin_Lin
Justin Long	http://en.wikipedia.org/wiki/Justin_Long
Justin Martyr	http://en.wikipedia.org/wiki/Justin_Martyr
Justin Rigali	http://en.wikipedia.org/wiki/Justin_Rigali
Justin Sane	http://en.wikipedia.org/wiki/Justin_Sane
Justin Theroux	http://en.wikipedia.org/wiki/Justin_Theroux
Justin Timberlake	http://en.wikipedia.org/wiki/Justin_Timberlake
Justin Tomlinson	http://en.wikipedia.org/wiki/Justin_Tomlinson
Justin Winsor	http://en.wikipedia.org/wiki/Justin_Winsor
Justine Bateman	http://en.wikipedia.org/wiki/Justine_Bateman
Justine Frischmann	http://en.wikipedia.org/wiki/Justine_Frischmann
Justine Greening	http://en.wikipedia.org/wiki/Justine_Greening
Justinian I	http://en.wikipedia.org/wiki/Justinian_I
Justo Jos� de Urquiza	http://en.wikipedia.org/wiki/Justo_Jos�_de_Urquiza
Justus Liebig	http://en.wikipedia.org/wiki/Justus_Liebig
Justus Lipsius	http://en.wikipedia.org/wiki/Justus_Lipsius
Justus Menius	http://en.wikipedia.org/wiki/Justus_Menius
K. Alex M�ller	http://en.wikipedia.org/wiki/K._Alex_Muller
K. Barry Sharpless	http://en.wikipedia.org/wiki/K._Barry_Sharpless
K. Eric Drexler	http://en.wikipedia.org/wiki/K._Eric_Drexler
K. R. Narayanan	http://en.wikipedia.org/wiki/K._R._Narayanan
K. T. Oslin	http://en.wikipedia.org/wiki/K._T._Oslin
K.D. Lang	http://en.wikipedia.org/wiki/K.d._lang
Kaavya Viswanathan	http://en.wikipedia.org/wiki/Kaavya_Viswanathan
Kadeem Hardison	http://en.wikipedia.org/wiki/Kadeem_Hardison
Kai Krause	http://en.wikipedia.org/wiki/Kai_Krause
Kai M. Siegbahn	http://en.wikipedia.org/wiki/Kai_M._Siegbahn
Kaiser Wilhelm	http://en.wikipedia.org/wiki/Wilhelm_II,_German_Emperor
Kak�	http://en.wikipedia.org/wiki/Kak�
Kal Penn	http://en.wikipedia.org/wiki/Kal_Penn
Kaley Cuoco	http://en.wikipedia.org/wiki/Kaley_Cuoco
Kalkot Mataskelekele	http://en.wikipedia.org/wiki/Kalkot_Mataskelekele
Kam Fong	http://en.wikipedia.org/wiki/Kam_Fong_Chun
Kamal Ahmed	http://en.wikipedia.org/wiki/Kamal_Ahmed
Kamal Al-Shennawi	http://en.wikipedia.org/wiki/Kamal_Al-Shennawi
Kamal Jumblatt	http://en.wikipedia.org/wiki/Kamal_Jumblatt
Kamal Nath	http://en.wikipedia.org/wiki/Kamal_Nath
Kamehameha I	http://en.wikipedia.org/wiki/Kamehameha_I
Kamla Persad-Bissessar	http://en.wikipedia.org/wiki/Kamla_Persad-Bissessar
Kane Hodder	http://en.wikipedia.org/wiki/Kane_Hodder
Kanye West	http://en.wikipedia.org/wiki/Kanye_West
Kareem Abdul-Jabbar	http://en.wikipedia.org/wiki/Kareem_Abdul-Jabbar
Karel Capek	http://en.wikipedia.org/wiki/Karel_%C4%8Capek
Karen Akers	http://en.wikipedia.org/wiki/Karen_Akers
Karen Allen	http://en.wikipedia.org/wiki/Karen_Allen
Karen Armstrong	http://en.wikipedia.org/wiki/Karen_Armstrong
Karen Black	http://en.wikipedia.org/wiki/Karen_Black
Karen Bradley	http://en.wikipedia.org/wiki/Karen_Bradley
Karen Buck	http://en.wikipedia.org/wiki/Karen_Buck
Karen Carpenter	http://en.wikipedia.org/wiki/Karen_Carpenter
Karen Czarnecki	http://en.wikipedia.org/wiki/Karen_Czarnecki
Karen Duffy	http://en.wikipedia.org/wiki/Karen_Duffy
Karen Finley	http://en.wikipedia.org/wiki/Karen_Finley
Karen Grassle	http://en.wikipedia.org/wiki/Karen_Grassle
Karen Hughes	http://en.wikipedia.org/wiki/Karen_Hughes
Karen Kilgariff	http://en.wikipedia.org/wiki/Karen_Kilgariff
Karen Lumley	http://en.wikipedia.org/wiki/Karen_Lumley
Karen Malina White	http://en.wikipedia.org/wiki/Karen_Malina_White
Karen Mantler	http://en.wikipedia.org/wiki/Karen_Mantler
Karen McCarthy	http://en.wikipedia.org/wiki/Karen_McCarthy
Karen Morley	http://en.wikipedia.org/wiki/Karen_Morley
Karen O	http://en.wikipedia.org/wiki/Karen_O
Karen Tumulty	http://en.wikipedia.org/wiki/Karen_Tumulty
Karen Valentine	http://en.wikipedia.org/wiki/Karen_Valentine
Karim Masimov	http://en.wikipedia.org/wiki/Karim_Masimov
Karina Lombard	http://en.wikipedia.org/wiki/Karina_Lombard
Karl Albrecht	http://en.wikipedia.org/wiki/Karl_Albrecht
Karl August von Hardenberg	http://en.wikipedia.org/wiki/Karl_August_von_Hardenberg
Karl Blake	http://en.wikipedia.org/wiki/Karl_Blake
Karl Carstens	http://en.wikipedia.org/wiki/Karl_Carstens
Karl Doenitz	http://en.wikipedia.org/wiki/Karl_Doenitz
Karl Ernst von Baer	http://en.wikipedia.org/wiki/Karl_Ernst_von_Baer
Karl Faberge	http://en.wikipedia.org/wiki/Karl_Faberge
Karl Gustav Jacobi	http://en.wikipedia.org/wiki/Karl_Gustav_Jacobi
Karl Lagerfeld	http://en.wikipedia.org/wiki/Karl_Lagerfeld
Karl Landsteiner	http://en.wikipedia.org/wiki/Karl_Landsteiner
Karl Malden	http://en.wikipedia.org/wiki/Karl_Malden
Karl Malone	http://en.wikipedia.org/wiki/Karl_Malone
Karl Mannheim	http://en.wikipedia.org/wiki/Karl_Mannheim
Karl Marx	http://en.wikipedia.org/wiki/Karl_Marx
Karl McCartney	http://en.wikipedia.org/wiki/Karl_McCartney
Karl Menninger	http://en.wikipedia.org/wiki/Karl_Menninger
Karl Philipp Moritz	http://en.wikipedia.org/wiki/Karl_Philipp_Moritz
Karl Popper	http://en.wikipedia.org/wiki/Karl_Popper
Karl Rove	http://en.wikipedia.org/wiki/Karl_Rove
Karl Shapiro	http://en.wikipedia.org/wiki/Karl_Shapiro
Karl Turner	http://en.wikipedia.org/wiki/Karl_Turner_(politician)
Karl Urban	http://en.wikipedia.org/wiki/Karl_Urban
Karl von Frisch	http://en.wikipedia.org/wiki/Karl_von_Frisch
Karl von Holtei	http://en.wikipedia.org/wiki/Karl_von_Holtei
Karl Ziegler	http://en.wikipedia.org/wiki/Karl_Ziegler
Karla Faye Tucker	http://en.wikipedia.org/wiki/Karla_Faye_Tucker
Karla Homolka	http://en.wikipedia.org/wiki/Karla_Homolka
Karl-Heinrich von Stuelpnagel	http://en.wikipedia.org/wiki/Karl-Heinrich_von_Stuelpnagel
Karlheinz Stockhausen	http://en.wikipedia.org/wiki/Karlheinz_Stockhausen
Karolina Kurkova	http://en.wikipedia.org/wiki/Karol%C3%ADna_Kurkov%C3%A1
Karpo Acimovic-Godina	http://en.wikipedia.org/wiki/Karpo_Acimovic-Godina
Kary Mullis	http://en.wikipedia.org/wiki/Kary_Mullis
Karyn Parsons	http://en.wikipedia.org/wiki/Karyn_Parsons
Kaspar Schwenkfeld	http://en.wikipedia.org/wiki/Kaspar_Schwenkfeld_von_Ossig
Katarina Witt	http://en.wikipedia.org/wiki/Katarina_Witt
Kate Ascher	http://en.wikipedia.org/wiki/Kate_Ascher
Kate Beckinsale	http://en.wikipedia.org/wiki/Kate_Beckinsale
Kate Bosworth	http://en.wikipedia.org/wiki/Kate_Bosworth
Kate Bush	http://en.wikipedia.org/wiki/Kate_Bush
Kate Capshaw	http://en.wikipedia.org/wiki/Kate_Capshaw
Kate Chopin	http://en.wikipedia.org/wiki/Kate_Chopin
Kate DiCamillo	http://en.wikipedia.org/wiki/Kate_DiCamillo
Kate Douglas Wiggin	http://en.wikipedia.org/wiki/Kate_Douglas_Wiggin
Kate Green	http://en.wikipedia.org/wiki/Kate_Green
Kate Greenaway	http://en.wikipedia.org/wiki/Kate_Greenaway
Kate Hoey	http://en.wikipedia.org/wiki/Kate_Hoey
Kate Hudson	http://en.wikipedia.org/wiki/Kate_Hudson 
Kate Jackson	http://en.wikipedia.org/wiki/Kate_Jackson
Kate Millett	http://en.wikipedia.org/wiki/Kate_Millett
Kate Moss	http://en.wikipedia.org/wiki/Kate_Moss
Kate Mulgrew	http://en.wikipedia.org/wiki/Kate_Mulgrew
Kate Nelligan	http://en.wikipedia.org/wiki/Kate_Nelligan
Kate O'Beirne	http://en.wikipedia.org/wiki/Kate_O%27Beirne
Kate O'Brien	http://en.wikipedia.org/wiki/Kate_O%27Brien
Kate Reid	http://en.wikipedia.org/wiki/Kate_Reid
Kate Smith	http://en.wikipedia.org/wiki/Kate_Smith
Kate Winslet	http://en.wikipedia.org/wiki/Kate_Winslet
Katey Sagal	http://en.wikipedia.org/wiki/Katey_Sagal
Katharine Anthony	http://en.wikipedia.org/wiki/Katharine_Anthony
Katharine Graham	http://en.wikipedia.org/wiki/Katharine_Graham
Katharine Hepburn	http://en.wikipedia.org/wiki/Katharine_Hepburn
Katharine Philips	http://en.wikipedia.org/wiki/Katharine_Philips
Katharine Ross	http://en.wikipedia.org/wiki/Katharine_Ross
Katharine Towne	http://en.wikipedia.org/wiki/Katharine_Towne
K�the Kollwitz	http://en.wikipedia.org/wiki/K%C3%A4the_Kollwitz
Katherine Anne Porter	http://en.wikipedia.org/wiki/Katherine_Anne_Porter
Katherine Dunham	http://en.wikipedia.org/wiki/Katherine_Dunham
Katherine Harris	http://en.wikipedia.org/wiki/Katherine_Harris
Katherine Heigl	http://en.wikipedia.org/wiki/Katherine_Heigl
Katherine Helmond	http://en.wikipedia.org/wiki/Katherine_Helmond
Katherine Kelly Lang	http://en.wikipedia.org/wiki/Katherine_Kelly_Lang
Katherine Lanpher	http://en.wikipedia.org/wiki/Katherine_Lanpher
Katherine Mansfield	http://en.wikipedia.org/wiki/Katherine_Mansfield
Katherine Moennig	http://en.wikipedia.org/wiki/Katherine_Moennig
Kathie Lee Gifford	http://en.wikipedia.org/wiki/Kathie_Lee_Gifford
Kathleen Beller	http://en.wikipedia.org/wiki/Kathleen_Beller
Kathleen Blanco	http://en.wikipedia.org/wiki/Kathleen_Blanco
Kathleen Hanna	http://en.wikipedia.org/wiki/Kathleen_Hanna
Kathleen Kennedy	http://en.wikipedia.org/wiki/Kathleen_Kennedy_%28film_producer%29
Kathleen Kennedy	http://en.wikipedia.org/wiki/Kathleen_Cavendish,_Marchioness_of_Hartington
Kathleen Q. Abernathy	http://en.wikipedia.org/wiki/Kathleen_Q._Abernathy
Kathleen Quinlan	http://en.wikipedia.org/wiki/Kathleen_Quinlan
Kathleen Sebelius	http://en.wikipedia.org/wiki/Kathleen_Sebelius
Kathleen Sullivan	http://en.wikipedia.org/wiki/Kathleen_Sullivan
Kathleen Turner	http://en.wikipedia.org/wiki/Kathleen_Turner
Kathleen Widdoes	http://en.wikipedia.org/wiki/Kathleen_Widdoes
Kathryn Bigelow	http://en.wikipedia.org/wiki/Kathryn_Bigelow
Kathryn Erbe	http://en.wikipedia.org/wiki/Kathryn_Erbe
Kathryn Grayson	http://en.wikipedia.org/wiki/Kathryn_Grayson
Kathryn Morris	http://en.wikipedia.org/wiki/Kathryn_Morris
Kathy Acker	http://en.wikipedia.org/wiki/Kathy_Acker
Kathy Baker	http://en.wikipedia.org/wiki/Kathy_Baker
Kathy Bates	http://en.wikipedia.org/wiki/Kathy_Bates
Kathy Castor	http://en.wikipedia.org/wiki/Kathy_Castor
Kathy Dahlkemper	http://en.wikipedia.org/wiki/Kathy_Dahlkemper 
Kathy Griffin	http://en.wikipedia.org/wiki/Kathy_Griffin
Kathy Ireland	http://en.wikipedia.org/wiki/Kathy_Ireland
Kathy Najimy	http://en.wikipedia.org/wiki/Kathy_Najimy
Kathy Valentine	http://en.wikipedia.org/wiki/Kathy_Valentine
Katie Cassidy	http://en.wikipedia.org/wiki/Katie_Cassidy
Katie Couric	http://en.wikipedia.org/wiki/Katie_Couric
Katie Holmes	http://en.wikipedia.org/wiki/Katie_Holmes
Katina Paxinou	http://en.wikipedia.org/wiki/Katina_Paxinou
Kato Kaelin	http://en.wikipedia.org/wiki/Kato_Kaelin
Katrina vanden Heuvel	http://en.wikipedia.org/wiki/Katrina_vanden_Heuvel
Katy Clark	http://en.wikipedia.org/wiki/Katy_Clark
Katy Jurado	http://en.wikipedia.org/wiki/Katy_Jurado
Kay Bailey Hutchison	http://en.wikipedia.org/wiki/Kay_Bailey_Hutchison
Kay Boyle	http://en.wikipedia.org/wiki/Kay_Boyle
Kay Francis	http://en.wikipedia.org/wiki/Kay_Francis
Kay Granger	http://en.wikipedia.org/wiki/Kay_Granger
Kay Hagan	http://en.wikipedia.org/wiki/Kay_Hagan
Kay Kendall	http://en.wikipedia.org/wiki/Kay_Kendall
Kay Kyser	http://en.wikipedia.org/wiki/Kay_Kyser
Kay Lenz	http://en.wikipedia.org/wiki/Kay_Lenz
Kay Nielsen	http://en.wikipedia.org/wiki/Kay_Nielsen
Kay Panabaker	http://en.wikipedia.org/wiki/Kay_Panabaker
Kay Walsh	http://en.wikipedia.org/wiki/Kay_Walsh
Kaye Ballard	http://en.wikipedia.org/wiki/Kaye_Ballard
Kaysone Phomvihane	http://en.wikipedia.org/wiki/Kaysone_Phomvihane
Kazimierz Marcinkiewicz	http://en.wikipedia.org/wiki/Kazimierz_Marcinkiewicz
Kazimir Malevich	http://en.wikipedia.org/wiki/Kazimir_Malevich
Kazuo Ishiguro	http://en.wikipedia.org/wiki/Kazuo_Ishiguro
Kazutoki Umezu	http://en.wikipedia.org/wiki/Kazutoki_Umezu
kd lang	http://en.wikipedia.org/wiki/kd_lang
Keanu Reeves	http://en.wikipedia.org/wiki/Keanu_Reeves
Keenan Wynn	http://en.wikipedia.org/wiki/Keenan_Wynn 
Keenen Ivory Wayans	http://en.wikipedia.org/wiki/Keenan_Ivory_Wayans
Keiichi Tsuchiya	http://en.wikipedia.org/wiki/Keiichi_Tsuchiya
Keir Dullea	http://en.wikipedia.org/wiki/Keir_Dullea
Keir Hardie	http://en.wikipedia.org/wiki/Keir_Hardie
Keira Knightley	http://en.wikipedia.org/wiki/Keira_Knightley
Keith Carradine	http://en.wikipedia.org/wiki/Keith_Carradine
Keith David	http://en.wikipedia.org/wiki/Keith_David
Keith Ellison	http://en.wikipedia.org/wiki/Keith_Ellison_%28politician%29
Keith Emerson	http://en.wikipedia.org/wiki/Keith_Emerson
Keith Fullerton Whitman	http://en.wikipedia.org/wiki/Keith_Fullerton_Whitman
Keith Haring	http://en.wikipedia.org/wiki/Keith_Haring
Keith Hernandez	http://en.wikipedia.org/wiki/Keith_Hernandez
Keith Knudsen	http://en.wikipedia.org/wiki/Keith_Knudsen
Keith Mitchell	http://en.wikipedia.org/wiki/Keith_Mitchell
Keith Moon	http://en.wikipedia.org/wiki/Keith_Moon
Keith Olbermann	http://en.wikipedia.org/wiki/Keith_Olbermann
Keith Richards	http://en.wikipedia.org/wiki/Keith_Richards
Keith Simpson	http://en.wikipedia.org/wiki/Keith_Simpson_%28politician%29
Keith Sweat	http://en.wikipedia.org/wiki/Keith_Sweat
Keith Urban	http://en.wikipedia.org/wiki/Keith_Urban
Keith Vaz	http://en.wikipedia.org/wiki/Keith_Vaz
Keith Waterhouse	http://en.wikipedia.org/wiki/Keith_Waterhouse
Keizo Obuchi	http://en.wikipedia.org/wiki/Keiz%C5%8D_Obuchi
Kel Mitchell	http://en.wikipedia.org/wiki/Kel_Mitchell
Kelley Deal	http://en.wikipedia.org/wiki/Kelley_Deal
Kelli White	http://en.wikipedia.org/wiki/Kelli_White
Kellie Martin	http://en.wikipedia.org/wiki/Kellie_Martin
Kellie Williams	http://en.wikipedia.org/wiki/Kellie_Williams
Ken Griffin	http://en.wikipedia.org/wiki/Kenneth_C._Griffin
Kenneth Burke	http://en.wikipedia.org/wiki/Kenneth_Burke
Kenneth Chenault	http://en.wikipedia.org/wiki/Kenneth_Chenault
Kenneth Clark	http://en.wikipedia.org/wiki/Kenneth_Clark
Kenneth Clarke	http://en.wikipedia.org/wiki/Kenneth_Clarke
Kenneth D. Lewis	http://en.wikipedia.org/wiki/Kenneth_D._Lewis
Kenneth E. Boulding	http://en.wikipedia.org/wiki/Kenneth_E._Boulding
Kenneth G. Wilson	http://en.wikipedia.org/wiki/Kenneth_G._Wilson
Kenneth Hall	http://en.wikipedia.org/wiki/Kenneth_O._Hall
Kenneth I	http://en.wikipedia.org/wiki/Kenneth_I
Kenneth I. Chenault	http://en.wikipedia.org/wiki/Kenneth_I._Chenault
Kenneth II	http://en.wikipedia.org/wiki/Kenneth_II_of_Scotland
Kenneth J. Arrow	http://en.wikipedia.org/wiki/Kenneth_J._Arrow
Kenneth J. Gray	http://en.wikipedia.org/wiki/Kenneth_J._Gray
Kenneth Kaunda	http://en.wikipedia.org/wiki/Kenneth_Kaunda
Kenneth Koch	http://en.wikipedia.org/wiki/Kenneth_Koch
Kenneth Mackenzie	http://en.wikipedia.org/wiki/Kenneth_%28Seaforth%29_Mackenzie
Kenneth More	http://en.wikipedia.org/wiki/Kenneth_More
Kenneth Parnell	http://en.wikipedia.org/wiki/Kenneth_Parnell
Kenneth Patchen	http://en.wikipedia.org/wiki/Kenneth_Patchen
Kenneth Rexroth	http://en.wikipedia.org/wiki/Kenneth_Rexroth
Kenneth Roberts	http://en.wikipedia.org/wiki/Kenneth_Roberts_%28author%29
Kenneth Tomlinson	http://en.wikipedia.org/wiki/Kenneth_Tomlinson
Kenneth Tynan	http://en.wikipedia.org/wiki/Kenneth_Tynan
Kenneth Williams	http://en.wikipedia.org/wiki/Kenneth_Williams
Kenny Anthony	http://en.wikipedia.org/wiki/Kenny_Anthony
Kenny Baker	http://en.wikipedia.org/wiki/Kenny_Baker
Kenny Chesney	http://en.wikipedia.org/wiki/Kenny_Chesney
Kenny Clarke	http://en.wikipedia.org/wiki/Kenny_Clarke
Kenny Dalglish	http://en.wikipedia.org/wiki/Kenny_Dalglish
Kenny G	http://en.wikipedia.org/wiki/Kenny_G
Kenny Guinn	http://en.wikipedia.org/wiki/Kenny_Guinn
Kenny Hickey	http://en.wikipedia.org/wiki/Kenny_Hickey
Kenny Hulshof	http://en.wikipedia.org/wiki/Kenny_Hulshof
Kenny Loggins	http://en.wikipedia.org/wiki/Kenny_Loggins
Kenny Lynch	http://en.wikipedia.org/wiki/Kenny_Lynch
Kenny Marchant	http://en.wikipedia.org/wiki/Kenny_Marchant
Kenny Rogers	http://en.wikipedia.org/wiki/Kenny_Rogers
Kenny Wayne Shepherd	http://en.wikipedia.org/wiki/Kenny_Wayne_Shepherd
Kent Conrad	http://en.wikipedia.org/wiki/Kent_Conrad
Kent Hovind	http://en.wikipedia.org/wiki/Kent_Hovind
Kent McCord	http://en.wikipedia.org/wiki/Kent_McCord
Kenyon Hopkins	http://en.wikipedia.org/wiki/Kenyon_Hopkins
Kenzaburo O�	http://en.wikipedia.org/wiki/Kenzabur%C5%8D_%C5%8Ce
Kenzo Tange	http://en.wikipedia.org/wiki/Kenzo_Tange
Keren Ann	http://en.wikipedia.org/wiki/Keren_Ann
Keri Russell	http://en.wikipedia.org/wiki/Keri_Russell
Kermit Roosevelt	http://en.wikipedia.org/wiki/Kermit_Roosevelt
Kerr Smith	http://en.wikipedia.org/wiki/Kerr_Smith
Kerri Kenney	http://en.wikipedia.org/wiki/Kerri_Kenney-Silver
Kerry King	http://en.wikipedia.org/wiki/Kerry_King
Kerry McCarthy	http://en.wikipedia.org/wiki/Kerry_McCarthy
Kerry Packer	http://en.wikipedia.org/wiki/Kerry_Packer
Kerry Washington	http://en.wikipedia.org/wiki/Kerry_Washington
Keshia Knight Pulliam	http://en.wikipedia.org/wiki/Keshia_Knight_Pulliam
Kessai Note	http://en.wikipedia.org/wiki/Kessai_Note
Kevan Jones	http://en.wikipedia.org/wiki/Kevan_Jones
Kevin Allison	http://en.wikipedia.org/wiki/Kevin_Allison
Kevin Ayers	http://en.wikipedia.org/wiki/Kevin_Ayers
Kevin Bacon	http://en.wikipedia.org/wiki/Kevin_Bacon
Kevin Barron	http://en.wikipedia.org/wiki/Kevin_Barron
Kevin Brady	http://en.wikipedia.org/wiki/Kevin_Brady
Kevin Brennan	http://en.wikipedia.org/wiki/Kevin_Brennan_%28politician%29
Kevin Connolly	http://en.wikipedia.org/wiki/Kevin_Connolly_%28actor%29
Kevin Cooper	http://en.wikipedia.org/wiki/Kevin_Cooper_%28inmate%29
Kevin Costner	http://en.wikipedia.org/wiki/Kevin_Costner
Kevin Dillon	http://en.wikipedia.org/wiki/Kevin_Dillon
Kevin Dobson	http://en.wikipedia.org/wiki/Kevin_Dobson
Kevin Eubanks	http://en.wikipedia.org/wiki/Kevin_Eubanks
Kevin Federline	http://en.wikipedia.org/wiki/Kevin_Federline
Kevin Garnett	http://en.wikipedia.org/wiki/Kevin_Garnett
Kevin Hagen	http://en.wikipedia.org/wiki/Kevin_Hagen
Kevin J. Anderson	http://en.wikipedia.org/wiki/Kevin_J._Anderson
Kevin J. Martin	http://en.wikipedia.org/wiki/Kevin_J._Martin
Kevin James	http://en.wikipedia.org/wiki/Kevin_James_%28actor%29
Kevin Keegan	http://en.wikipedia.org/wiki/Kevin_Keegan
Kevin Kline	http://en.wikipedia.org/wiki/Kevin_Kline
Kevin McCarthy	http://en.wikipedia.org/wiki/Kevin_McCarthy_%28actor%29
Kevin McCarthy	http://en.wikipedia.org/wiki/Kevin_McCarthy_%28California%29
Kevin McDonald	http://en.wikipedia.org/wiki/Kevin_McDonald
Kevin Mitnick	http://en.wikipedia.org/wiki/Kevin_Mitnick
Kevin Nealon	http://en.wikipedia.org/wiki/Kevin_Nealon
Kevin Peter Hall	http://en.wikipedia.org/wiki/Kevin_Peter_Hall
Kevin Phillips	http://en.wikipedia.org/wiki/Kevin_Phillips_%28political_commentator%29
Kevin Pollak	http://en.wikipedia.org/wiki/Kevin_Pollak
Kevin Poulsen	http://en.wikipedia.org/wiki/Kevin_Poulsen
Kevin Richardson	http://en.wikipedia.org/wiki/Kevin_Richardson_%28musician%29
Kevin Rollins	http://en.wikipedia.org/wiki/Kevin_Rollins
Kevin Rudd	http://en.wikipedia.org/wiki/Kevin_Rudd
Kevin Shelley	http://en.wikipedia.org/wiki/Kevin_Shelley
Kevin Shields	http://en.wikipedia.org/wiki/Kevin_Shields
Kevin Smith	http://en.wikipedia.org/wiki/Kevin_Smith
Kevin Sorbo	http://en.wikipedia.org/wiki/Kevin_Sorbo
Kevin Spacey	http://en.wikipedia.org/wiki/Kevin_Spacey
Kevin Trudeau	http://en.wikipedia.org/wiki/Kevin_Trudeau
Kevin W. Sharer	http://en.wikipedia.org/wiki/Kevin_W._Sharer
Kevin Williamson	http://en.wikipedia.org/wiki/Kevin_Williamson_%28screenwriter%29
Kevin Zegers	http://en.wikipedia.org/wiki/Kevin_Zegers
Keyshia Cole	http://en.wikipedia.org/wiki/Keyshia_Cole
Khaled Mashaal	http://en.wikipedia.org/wiki/Khaled_Mashaal
Khaleda Zia	http://en.wikipedia.org/wiki/Khaleda_Zia
Khalid Mahmood	http://en.wikipedia.org/wiki/Khalid_Mahmood
Khalid Shaikh Mohammed	http://en.wikipedia.org/wiki/Khalid_Shaikh_Mohammed
Khalifa ibn Salman Ali Khalifa	http://en.wikipedia.org/wiki/Khalifah_ibn_Sulman_Al_Khalifah
Khalifa ibn Zayed Al Nahayan	http://en.wikipedia.org/wiki/Khalifa_ibn_Zayed_al-Nahayan
Khalil Gibran	http://en.wikipedia.org/wiki/Khalil_Gibran
Khamtai Siphandon	http://en.wikipedia.org/wiki/Khamtai_Siphandon
Khandi Alexander	http://en.wikipedia.org/wiki/Khandi_Alexander
Khigh Dhiegh	http://en.wikipedia.org/wiki/Khigh_Dhiegh
Kid 606	http://en.wikipedia.org/wiki/Kid_606
Kid Koala	http://en.wikipedia.org/wiki/Kid_Koala
Kid Loco	http://en.wikipedia.org/wiki/Kid_Loco
Kid Rock	http://en.wikipedia.org/wiki/Kid_Rock
Kiefer Sutherland	http://en.wikipedia.org/wiki/Kiefer_Sutherland
Kieran Culkin	http://en.wikipedia.org/wiki/Kieran_Culkin
Kieran Hebden	http://en.wikipedia.org/wiki/Kieran_Hebden
Kiichi Miyazawa	http://en.wikipedia.org/wiki/Kiichi_Miyazawa
Kika de la Garza	http://en.wikipedia.org/wiki/Kika_de_la_Garza
Killer Kowalski	http://en.wikipedia.org/wiki/Killer_Kowalski
Killer Mike	http://en.wikipedia.org/wiki/Killer_Mike
Kim Alexis	http://en.wikipedia.org/wiki/Kim_Alexis
Kim Basinger	http://en.wikipedia.org/wiki/Kim_Basinger
Kim Campbell	http://en.wikipedia.org/wiki/Kim_Campbell
Kim Carnes	http://en.wikipedia.org/wiki/Kim_Carnes
Kim Cattrall	http://en.wikipedia.org/wiki/Kim_Cattrall
Kim Dae-Jung	http://en.wikipedia.org/wiki/Kim_Dae-jung
Kim Darby	http://en.wikipedia.org/wiki/Kim_Darby
Kim Deal	http://en.wikipedia.org/wiki/Kim_Deal
Kim Delaney	http://en.wikipedia.org/wiki/Kim_Delaney
Kim Fields	http://en.wikipedia.org/wiki/Kim_Fields
Kim Gordon	http://en.wikipedia.org/wiki/Kim_Gordon
Kim Hunter	http://en.wikipedia.org/wiki/Kim_Hunter
Kim Il Sung	http://en.wikipedia.org/wiki/Kim_Il-sung
Kim Jong Il	http://en.wikipedia.org/wiki/Kim_Jong-il
Kim Novak	http://en.wikipedia.org/wiki/Kim_Novak
Kim Peek	http://en.wikipedia.org/wiki/Kim_Peek
Kim Philby	http://en.wikipedia.org/wiki/Kim_Philby
Kim Richards	http://en.wikipedia.org/wiki/Kim_Richards
Kim Weston	http://en.wikipedia.org/wiki/Kim_Weston
Kim Wilde	http://en.wikipedia.org/wiki/Kim_Wilde
Kim Yong-nam	http://en.wikipedia.org/wiki/Kim_Yong-nam
Kim Young Sam	http://en.wikipedia.org/wiki/Kim_Young-sam
Kim Zimmer	http://en.wikipedia.org/wiki/Kim_Zimmer
Kimberley Rew	http://en.wikipedia.org/wiki/Kimberley_Rew
Kimberly Dozier	http://en.wikipedia.org/wiki/Kimberly_Dozier
Kimberly Elise	http://en.wikipedia.org/wiki/Kimberly_Elise
Kimberly Williams	http://en.wikipedia.org/wiki/Kimberly_Williams-Paisley
Kimi Raikkonen	http://en.wikipedia.org/wiki/Kimi_R%C3%A4ikk%C3%B6nen
Kimora Lee Simmons	http://en.wikipedia.org/wiki/Kimora_Lee_Simmons
Kin Hubbard	http://en.wikipedia.org/wiki/Kin_Hubbard
King Abdullah	http://en.wikipedia.org/wiki/Abdullah_of_Saudi_Arabia
King Abdullah II	http://en.wikipedia.org/wiki/King_Abdullah_II
King Ad-Rock	http://en.wikipedia.org/wiki/King_Ad-Rock
King Albert II	http://en.wikipedia.org/wiki/Albert_II_of_Belgium
King Alfred the Great	http://en.wikipedia.org/wiki/Alfred_the_Great
King Athelstan	http://en.wikipedia.org/wiki/King_Athelstan
King Canute	http://en.wikipedia.org/wiki/King_Canute
King Carl XVI Gustaf	http://en.wikipedia.org/wiki/King_Carl_XVI_Gustaf
King Charles I	http://en.wikipedia.org/wiki/Charles_I_of_England
King Charles II	http://en.wikipedia.org/wiki/Charles_II_of_England
King Charles XII	http://en.wikipedia.org/wiki/Charles_XII_of_Sweden
King Diamond	http://en.wikipedia.org/wiki/King_Diamond
King Donovan	http://en.wikipedia.org/wiki/King_Donovan
King Edgar I	http://en.wikipedia.org/wiki/King_Edgar
King Edmund I	http://en.wikipedia.org/wiki/Edmund_I_of_England
King Edmund II	http://en.wikipedia.org/wiki/Edmund_II
King Edred	http://en.wikipedia.org/wiki/Eadred_of_England
King Edward I	http://en.wikipedia.org/wiki/Edward_I_of_England
King Edward II	http://en.wikipedia.org/wiki/Edward_II_of_England
King Edward III	http://en.wikipedia.org/wiki/Edward_III_of_England
King Edward IV	http://en.wikipedia.org/wiki/Edward_IV_of_England
King Edward the Elder	http://en.wikipedia.org/wiki/Edward_the_Elder
King Edward V	http://en.wikipedia.org/wiki/Edward_V_of_England
King Edward VI	http://en.wikipedia.org/wiki/Edward_VI_of_England
King Edward VII	http://en.wikipedia.org/wiki/Edward_VII_of_the_United_Kingdom
King Edward VIII	http://en.wikipedia.org/wiki/Edward_VIII_of_the_United_Kingdom
King Edwy	http://en.wikipedia.org/wiki/Eadwig_of_England
King Ethelred II	http://en.wikipedia.org/wiki/Ethelred_II
King Ethelweard	http://en.wikipedia.org/wiki/%C3%86lfweard_of_Wessex
King Fahd	http://en.wikipedia.org/wiki/King_Fahd
King Ferdinand II	http://en.wikipedia.org/wiki/Ferdinand_II_of_Aragon
King Frederick I	http://en.wikipedia.org/wiki/Frederick_I,_Holy_Roman_Emperor
King George I	http://en.wikipedia.org/wiki/George_I_of_Great_Britain
King George II	http://en.wikipedia.org/wiki/George_II_of_Great_Britain
King George III	http://en.wikipedia.org/wiki/George_III_of_the_United_Kingdom
King George IV	http://en.wikipedia.org/wiki/George_IV_of_the_United_Kingdom
King George Tupou V	http://en.wikipedia.org/wiki/George_Tupou_V
King George V	http://en.wikipedia.org/wiki/George_V_of_the_United_Kingdom
King George VI	http://en.wikipedia.org/wiki/George_VI_of_the_United_Kingdom
King Gyanendra	http://en.wikipedia.org/wiki/Gyanendra_of_Nepal
King Harald V	http://en.wikipedia.org/wiki/Harald_V_of_Norway
King Harold II	http://en.wikipedia.org/wiki/Harold_Godwinson
King Harthacnut	http://en.wikipedia.org/wiki/Harthacnut_%281020%E2%80%931042%29
King Henry I	http://en.wikipedia.org/wiki/Henry_I_of_England
King Henry II	http://en.wikipedia.org/wiki/Henry_II_of_England
King Henry III	http://en.wikipedia.org/wiki/Henry_III_of_England
King Henry IV	http://en.wikipedia.org/wiki/Henry_IV_of_England
King Henry V	http://en.wikipedia.org/wiki/Henry_V_of_England
King Henry VI	http://en.wikipedia.org/wiki/Henry_VI_of_England
King Henry VII	http://en.wikipedia.org/wiki/Henry_VII_of_England
King Henry VIII	http://en.wikipedia.org/wiki/Henry_VIII_of_England
King Hussein I	http://en.wikipedia.org/wiki/Hussein_I
King James I	http://en.wikipedia.org/wiki/James_I_of_England
King James II	http://en.wikipedia.org/wiki/James_II_of_England
King John Lackland	http://en.wikipedia.org/wiki/John_of_England
King Juan Carlos I	http://en.wikipedia.org/wiki/Juan_Carlos_I_of_Spain
King Letsie III	http://en.wikipedia.org/wiki/Letsie_III_of_Lesotho
King Mohammed VI	http://en.wikipedia.org/wiki/Mohammed_VI_of_Morocco
King Mswati III	http://en.wikipedia.org/wiki/Mswati_III_of_Swaziland
King Richard II	http://en.wikipedia.org/wiki/Richard_II_of_England
King Richard III	http://en.wikipedia.org/wiki/Richard_III_of_England
King Richard the Lionheart	http://en.wikipedia.org/wiki/Richard_the_Lionheart
King Stephen	http://en.wikipedia.org/wiki/King_Stephen_of_England
King Sunny Ade	http://en.wikipedia.org/wiki/King_Sunny_Ad%C3%A9
King Vidor	http://en.wikipedia.org/wiki/King_Vidor
King William II	http://en.wikipedia.org/wiki/William_II_of_England
King William IV	http://en.wikipedia.org/wiki/William_IV_of_the_United_Kingdom
Kingsley Amis	http://en.wikipedia.org/wiki/Kingsley_Amis
Kinky Friedman	http://en.wikipedia.org/wiki/Kinky_Friedman
Kinya Aikawa	http://en.wikipedia.org/wiki/Kinya_Aikawa
Kip Pardue	http://en.wikipedia.org/wiki/Kip_Pardue
Kip Winger	http://en.wikipedia.org/wiki/Kip_Winger
Kira Roessler	http://en.wikipedia.org/wiki/Kira_Roessler
Kirby Puckett	http://en.wikipedia.org/wiki/Kirby_Puckett
Kirk Acevedo	http://en.wikipedia.org/wiki/Kirk_Acevedo
Kirk Alyn	http://en.wikipedia.org/wiki/Kirk_Alyn
Kirk Cameron	http://en.wikipedia.org/wiki/Kirk_Cameron
Kirk Douglas	http://en.wikipedia.org/wiki/Kirk_Douglas
Kirk Fordice	http://en.wikipedia.org/wiki/Kirk_Fordice
Kirk Franklin	http://en.wikipedia.org/wiki/Kirk_Franklin
Kirk Gibson	http://en.wikipedia.org/wiki/Kirk_Gibson
Kirk Hammett	http://en.wikipedia.org/wiki/Kirk_Hammett
Kirk Kerkorian	http://en.wikipedia.org/wiki/Kirk_Kerkorian
Kirsten Dunst	http://en.wikipedia.org/wiki/Kirsten_Dunst
Kirsten Gillibrand	http://en.wikipedia.org/wiki/Kirsten_Gillibrand
Kirsten Storms	http://en.wikipedia.org/wiki/Kirsten_Storms
Kirstie Alley	http://en.wikipedia.org/wiki/Kirstie_Alley
Kit Bond	http://en.wikipedia.org/wiki/Kit_Bond
Kit Carson	http://en.wikipedia.org/wiki/Kit_Carson
Kit Clayton	http://en.wikipedia.org/wiki/Kit_Clayton
Kitty Carlisle	http://en.wikipedia.org/wiki/Kitty_Carlisle
Kitty Dukakis	http://en.wikipedia.org/wiki/Kitty_Dukakis
Kitty Genovese	http://en.wikipedia.org/wiki/Kitty_Genovese
Kitty Kelley	http://en.wikipedia.org/wiki/Kitty_Kelley
Kitty Wells	http://en.wikipedia.org/wiki/Kitty_Wells
Kjell Magne Bondevik	http://en.wikipedia.org/wiki/Kjell_Magne_Bondevik
Klas Pontus Arnoldson	http://en.wikipedia.org/wiki/Klas_Pontus_Arnoldson
Klaus Barbie	http://en.wikipedia.org/wiki/Klaus_Barbie
Klaus Fuchs	http://en.wikipedia.org/wiki/Klaus_Fuchs
Klaus Kinkel	http://en.wikipedia.org/wiki/Klaus_Kinkel
Klaus Kinski	http://en.wikipedia.org/wiki/Klaus_Kinski
Klaus Nomi	http://en.wikipedia.org/wiki/Klaus_Nomi
Klaus Schulze	http://en.wikipedia.org/wiki/Klaus_Schulze
Klaus Tsch�tscher	http://en.wikipedia.org/wiki/Klaus_Tsch%C3%Bctscher
Klaus von Klitzing	http://en.wikipedia.org/wiki/Klaus_von_Klitzing
Klemens Wenzel von Metternich	http://en.wikipedia.org/wiki/Klemens_Wenzel_von_Metternich
Knut Hamsun	http://en.wikipedia.org/wiki/Knut_Hamsun
Knute Rockne	http://en.wikipedia.org/wiki/Knute_Rockne
Kobe Bryant	http://en.wikipedia.org/wiki/Kobe_Bryant
Kofi Annan	http://en.wikipedia.org/wiki/Kofi_Annan
Kofi Awoonor	http://en.wikipedia.org/wiki/Kofi_Awoonor
Koichi Tanaka	http://en.wikipedia.org/wiki/Koichi_Tanaka
Kon Artis	http://en.wikipedia.org/wiki/Kon_Artis
Konrad Adenauer	http://en.wikipedia.org/wiki/Konrad_Adenauer
Konrad Lorenz	http://en.wikipedia.org/wiki/Konrad_Lorenz
Konrad Mutian	http://en.wikipedia.org/wiki/Konrad_Mutian
Konrad von Gesner	http://en.wikipedia.org/wiki/Konrad_von_Gesner
Konstantin Chernenko	http://en.wikipedia.org/wiki/Konstantin_Chernenko
Konstantin E. Tsiolkovsky	http://en.wikipedia.org/wiki/Konstantin_E._Tsiolkovsky
Konstantin Fehrenbach	http://en.wikipedia.org/wiki/Konstantin_Fehrenbach
Konstantin von Neurath	http://en.wikipedia.org/wiki/Konstantin_von_Neurath
Kool G Rap	http://en.wikipedia.org/wiki/Kool_G_Rap
Kool Keith	http://en.wikipedia.org/wiki/Kool_Keith
Kool Moe Dee	http://en.wikipedia.org/wiki/Kool_Moe_Dee
Kordell Stewart	http://en.wikipedia.org/wiki/Kordell_Stewart
Korhan Abay	http://en.wikipedia.org/wiki/Korhan_Abay
Koumei Nakamura	http://en.wikipedia.org/wiki/Koumei_Nakamura
Kris Hopkins	http://en.wikipedia.org/wiki/Kris_Hopkins
Kris Kristofferson	http://en.wikipedia.org/wiki/Kris_Kristofferson
Krist Novoselic	http://en.wikipedia.org/wiki/Krist_Novoselic
Krista Allen	http://en.wikipedia.org/wiki/Krista_Allen
Kristanna Loken	http://en.wikipedia.org/wiki/Kristanna_Loken
Kristeen Young	http://en.wikipedia.org/wiki/Kristeen_Young
Kristen Bell	http://en.wikipedia.org/wiki/Kristen_Bell
Kristen Johnston	http://en.wikipedia.org/wiki/Kristen_Johnston
Kristen Pfaff	http://en.wikipedia.org/wiki/Kristen_Pfaff
Kristi Yamaguchi	http://en.wikipedia.org/wiki/Kristi_Yamaguchi
Kristian Alfonso	http://en.wikipedia.org/wiki/Kristian_Alfonso
Kristin Chenoweth	http://en.wikipedia.org/wiki/Kristin_Chenoweth
Kristin Davis	http://en.wikipedia.org/wiki/Kristin_Davis
Kristin Hersh	http://en.wikipedia.org/wiki/Kristin_Hersh
Kristin Kreuk	http://en.wikipedia.org/wiki/Kristin_Kreuk
Kristin Lehman	http://en.wikipedia.org/wiki/Kristin_Lehman
Kristin Scott Thomas	http://en.wikipedia.org/wiki/Kristin_Scott_Thomas
Kristina Adolphson	http://en.wikipedia.org/wiki/Kristina_Adolphson
Kristina Wagner	http://en.wikipedia.org/wiki/Kristina_Wagner
Kristine Kathryn Rusch	http://en.wikipedia.org/wiki/Kristine_Kathryn_Rusch
Kristy McNichol	http://en.wikipedia.org/wiki/Kristy_McNichol
Kristy Swanson	http://en.wikipedia.org/wiki/Kristy_Swanson
Krzysztof Penderecki	http://en.wikipedia.org/wiki/Krzysztof_Penderecki
Kublai Khan	http://en.wikipedia.org/wiki/Kublai_Khan
Kumar Sangakkara	http://en.wikipedia.org/wiki/Kumar_Sangakkara
Kurmanbek Bakiyev	http://en.wikipedia.org/wiki/Kurmanbek_Bakiyev
Kurt Alder	http://en.wikipedia.org/wiki/Kurt_Alder
Kurt Angle	http://en.wikipedia.org/wiki/Kurt_Angle
Kurt Cobain	http://en.wikipedia.org/wiki/Kurt_Cobain
Kurt Eichenwald	http://en.wikipedia.org/wiki/Kurt_Eichenwald
Kurt Georg Kiesinger	http://en.wikipedia.org/wiki/Kurt_Georg_Kiesinger
Kurt G�del	http://en.wikipedia.org/wiki/Kurt_G%C3%B6del
Kurt Loder	http://en.wikipedia.org/wiki/Kurt_Loder
Kurt Nilsen	http://en.wikipedia.org/wiki/Kurt_Nilsen
Kurt Russell	http://en.wikipedia.org/wiki/Kurt_Russell
Kurt Schrader	http://en.wikipedia.org/wiki/Kurt_Schrader
Kurt Schwitters	http://en.wikipedia.org/wiki/Kurt_Schwitters
Kurt Student	http://en.wikipedia.org/wiki/Kurt_Student
Kurt von Schleicher	http://en.wikipedia.org/wiki/Kurt_von_Schleicher
Kurt Vonnegut	http://en.wikipedia.org/wiki/Kurt_Vonnegut
Kurt Wüthrich	http://en.wikipedia.org/wiki/Kurt_W%C3%BCthrich
Kurt Waldheim	http://en.wikipedia.org/wiki/Kurt_Waldheim
Kurt Weill	http://en.wikipedia.org/wiki/Kurt_Weill
Kurtis Blow	http://en.wikipedia.org/wiki/Kurtis_Blow
Kurtwood Smith	http://en.wikipedia.org/wiki/Kurtwood_Smith
Kwame Anthony Appiah	http://en.wikipedia.org/wiki/Kwame_Anthony_Appiah
Kwame Nkrumah	http://en.wikipedia.org/wiki/Kwame_Nkrumah
Kwasi Kwarteng	http://en.wikipedia.org/wiki/Kwasi_Kwarteng
Kweisi Mfume	http://en.wikipedia.org/wiki/Kweisi_Mfume
Kyan Douglas	http://en.wikipedia.org/wiki/Kyan_Douglas
Kyla Pratt	http://en.wikipedia.org/wiki/Kyla_Pratt
Kyle Boller	http://en.wikipedia.org/wiki/Kyle_Boller
Kyle Chandler	http://en.wikipedia.org/wiki/Kyle_Chandler
Kyle Gass	http://en.wikipedia.org/wiki/Kyle_Gass
Kyle MacLachlan	http://en.wikipedia.org/wiki/Kyle_MacLachlan
Kyle Massey	http://en.wikipedia.org/wiki/Kyle_Massey
Kyle Secor	http://en.wikipedia.org/wiki/Kyle_Secor
Kylie Minogue	http://en.wikipedia.org/wiki/Kylie_Minogue
Kyra Sedgwick	http://en.wikipedia.org/wiki/Kyra_Sedgwick
L. Douglas Wilder	http://en.wikipedia.org/wiki/L._Douglas_Wilder
L. Frank Baum	http://en.wikipedia.org/wiki/L._Frank_Baum
L. Lowry Mays	http://en.wikipedia.org/wiki/L._Lowry_Mays
L. P. Hartley	http://en.wikipedia.org/wiki/L._P._Hartley
L. Patrick Gray	http://en.wikipedia.org/wiki/L._Patrick_Gray
L. Paul Bremer	http://en.wikipedia.org/wiki/L._Paul_Bremer
L. Ron Hubbard	http://en.wikipedia.org/wiki/L._Ron_Hubbard
L. Sprague de Camp	http://en.wikipedia.org/wiki/L._Sprague_de_Camp
La Monte Young	http://en.wikipedia.org/wiki/La_Monte_Young
La Toya Jackson	http://en.wikipedia.org/wiki/La_Toya_Jackson
La Voisin	http://en.wikipedia.org/wiki/La_Voisin
Lacey Chabert	http://en.wikipedia.org/wiki/Lacey_Chabert
Laci Peterson	http://en.wikipedia.org/wiki/Laci_Peterson
Lacy Clay	http://en.wikipedia.org/wiki/Lacy_Clay
Lacy J. Dalton	http://en.wikipedia.org/wiki/Lacy_J._Dalton
Ladislas I	http://en.wikipedia.org/wiki/Ladislas_I_of_Hungary
Ladislas IV	http://en.wikipedia.org/wiki/Ladislas_IV
Ladislas V	http://en.wikipedia.org/wiki/Ladislas_V
Ladislav Kl�ma	http://en.wikipedia.org/wiki/Ladislav_Kl%C3%Adma
Lady Bird Johnson	http://en.wikipedia.org/wiki/Lady_Bird_Johnson
Lady Diana	http://en.wikipedia.org/wiki/Lady_Diana
Lady Gaga	http://en.wikipedia.org/wiki/Lady_Gaga
Lady Jane Grey	http://en.wikipedia.org/wiki/Lady_Jane_Grey
Lady Mary Wortley Montagu	http://en.wikipedia.org/wiki/Lady_Mary_Wortley_Montagu
Lady Saw	http://en.wikipedia.org/wiki/Lady_Saw
Laetitia Casta	http://en.wikipedia.org/wiki/Laetitia_Casta
Laetitia Sadier	http://en.wikipedia.org/wiki/Laetitia_Sadier
Lafcadio Hearn	http://en.wikipedia.org/wiki/Lafcadio_Hearn
Laffit Pincay	http://en.wikipedia.org/wiki/Laffit_Pincay,_Jr.
Laisenia Qarase	http://en.wikipedia.org/wiki/Laisenia_Qarase
Lakhdar Brahimi	http://en.wikipedia.org/wiki/Lakhdar_Brahimi
Lakshmi Mittal	http://en.wikipedia.org/wiki/Lakshmi_Mittal
Lalla Ward	http://en.wikipedia.org/wiki/Lalla_Ward
Lally Weymouth	http://en.wikipedia.org/wiki/Lally_Weymouth
Lamar Alexander	http://en.wikipedia.org/wiki/Lamar_Alexander
Lamar Hunt	http://en.wikipedia.org/wiki/Lamar_Hunt
Lamar Smith	http://en.wikipedia.org/wiki/Lamar_S._Smith
Lamb Gaede	http://en.wikipedia.org/wiki/Lamb_Gaede
Lamont Bentley	http://en.wikipedia.org/wiki/Lamont_Bentley
Lana Turner	http://en.wikipedia.org/wiki/Lana_Turner
Lana Wood	http://en.wikipedia.org/wiki/Lana_Wood
Lance Acord	http://en.wikipedia.org/wiki/Lance_Acord
Lance Armstrong	http://en.wikipedia.org/wiki/Lance_Armstrong
Lance Bass	http://en.wikipedia.org/wiki/Lance_Bass
Lance Burton	http://en.wikipedia.org/wiki/Lance_Burton
Lance Henriksen	http://en.wikipedia.org/wiki/Lance_Henriksen
Lance Ito	http://en.wikipedia.org/wiki/Lance_Ito
Lance Kerwin	http://en.wikipedia.org/wiki/Lance_Kerwin
Lance Reddick	http://en.wikipedia.org/wiki/Lance_Reddick
Lance Rentzel	http://en.wikipedia.org/wiki/Lance_Rentzel
Landon Parvin	http://en.wikipedia.org/wiki/Landon_Parvin
Lane Evans	http://en.wikipedia.org/wiki/Lane_Evans
Lane Kirkland	http://en.wikipedia.org/wiki/Lane_Kirkland
Lane Smith	http://en.wikipedia.org/wiki/Lane_Smith
Lanford Wilson	http://en.wikipedia.org/wiki/Lanford_Wilson
Langston Hughes	http://en.wikipedia.org/wiki/Langston_Hughes
Lani Guinier	http://en.wikipedia.org/wiki/Lani_Guinier
Lani Hall	http://en.wikipedia.org/wiki/Lani_Hall
Lansana Cont�	http://en.wikipedia.org/wiki/Lansana_Cont%C3%A9
Lara Flynn Boyle	http://en.wikipedia.org/wiki/Lara_Flynn_Boyle
Lara Logan	http://en.wikipedia.org/wiki/Lara_Logan
Laraine Day	http://en.wikipedia.org/wiki/Laraine_Day
Laraine Newman	http://en.wikipedia.org/wiki/Laraine_Newman
Larenz Tate	http://en.wikipedia.org/wiki/Larenz_Tate
Larisa Oleynik	http://en.wikipedia.org/wiki/Larisa_Oleynik
Lark Voorhies	http://en.wikipedia.org/wiki/Lark_Voorhies
Larry A. Thompson	http://en.wikipedia.org/wiki/Larry_A._Thompson
Larry Adler	http://en.wikipedia.org/wiki/Larry_Adler
Larry Bird	http://en.wikipedia.org/wiki/Larry_Bird
Larry Bossidy	http://en.wikipedia.org/wiki/Larry_Bossidy
Larry Buchanan	http://en.wikipedia.org/wiki/Larry_Buchanan
Larry Collins	http://en.wikipedia.org/wiki/Larry_Collins_%28writer%29
Larry Combest	http://en.wikipedia.org/wiki/Larry_Combest
Larry Craig	http://en.wikipedia.org/wiki/Larry_Craig
Larry Csonka	http://en.wikipedia.org/wiki/Larry_Csonka
Larry David	http://en.wikipedia.org/wiki/Larry_David
Larry Elder	http://en.wikipedia.org/wiki/Larry_Elder
Larry Ellison	http://en.wikipedia.org/wiki/Larry_Ellison
Larry Fine	http://en.wikipedia.org/wiki/Larry_Fine
Larry Flynt	http://en.wikipedia.org/wiki/Larry_Flynt
Larry Fortensky	http://en.wikipedia.org/wiki/Larry_Fortensky
Larry Gatlin	http://en.wikipedia.org/wiki/Larry_Gatlin
Larry Gelbart	http://en.wikipedia.org/wiki/Larry_Gelbart
Larry Graham	http://en.wikipedia.org/wiki/Larry_Graham
Larry Hagman	http://en.wikipedia.org/wiki/Larry_Hagman
Larry Harvey	http://en.wikipedia.org/wiki/Larry_Harvey
Larry Holmes	http://en.wikipedia.org/wiki/Larry_Holmes
Larry Hovis	http://en.wikipedia.org/wiki/Larry_Hovis
Larry J. Hopkins	http://en.wikipedia.org/wiki/Larry_J._Hopkins
Larry King	http://en.wikipedia.org/wiki/Larry_King
Larry Kissell	http://en.wikipedia.org/wiki/Larry_Kissell
Larry Lea	http://en.wikipedia.org/wiki/Larry_Lea
Larry Levan	http://en.wikipedia.org/wiki/Larry_Levan
Larry Lindsey	http://en.wikipedia.org/wiki/Larry_Lindsey
Larry Linville	http://en.wikipedia.org/wiki/Larry_Linville
Larry Manetti	http://en.wikipedia.org/wiki/Larry_Manetti
Larry Mantle	http://en.wikipedia.org/wiki/Larry_Mantle
Larry McMurtry	http://en.wikipedia.org/wiki/Larry_McMurtry
Larry Miller	http://en.wikipedia.org/wiki/Larry_Miller_%28actor%29
Larry Mullen	http://en.wikipedia.org/wiki/Larry_Mullen,_Jr.
Larry Niven	http://en.wikipedia.org/wiki/Larry_Niven
Larry Norman	http://en.wikipedia.org/wiki/Larry_Norman
Larry Page	http://en.wikipedia.org/wiki/Larry_Page
Larry Parks	http://en.wikipedia.org/wiki/Larry_Parks
Larry Peerce	http://en.wikipedia.org/wiki/Larry_Peerce
Larry Pressler	http://en.wikipedia.org/wiki/Larry_Pressler
Larry Roberts	http://en.wikipedia.org/wiki/Lawrence_Roberts_%28scientist%29
Larry Speakes	http://en.wikipedia.org/wiki/Larry_Speakes
Larry Storch	http://en.wikipedia.org/wiki/Larry_Storch
Larry The Cable Guy	http://en.wikipedia.org/wiki/Larry_the_Cable_Guy
Larry Wachowski	http://en.wikipedia.org/wiki/Larry_Wachowski
Larry Wall	http://en.wikipedia.org/wiki/Larry_Wall
Larry Wilcox	http://en.wikipedia.org/wiki/Larry_Wilcox
Larry Wilkerson	http://en.wikipedia.org/wiki/Larry_Wilkerson
Larry Williams	http://en.wikipedia.org/wiki/Larry_Williams
Larry Woiwode	http://en.wikipedia.org/wiki/Larry_Woiwode
Lars Frederiksen	http://en.wikipedia.org/wiki/Lars_Frederiksen
Lars L�kke Rasmussen	http://en.wikipedia.org/wiki/Lars_L%C3%B8kke_Rasmussen
Lars Onsager	http://en.wikipedia.org/wiki/Lars_Onsager
Lars Ulrich	http://en.wikipedia.org/wiki/Lars_Ulrich
Lars von Trier	http://en.wikipedia.org/wiki/Lars_von_Trier
Lasse Braun	http://en.wikipedia.org/wiki/Lasse_Braun
Lasse Hallstrom	http://en.wikipedia.org/wiki/Lasse_Hallstr%C3%B6m
L�szl� Moholy-Nagy	http://en.wikipedia.org/wiki/L%e1szl%f3_Moholy-Nagy
L�szl� S�lyom	http://en.wikipedia.org/wiki/L%e1szl%f3_S%f3lyom
LaToya London	http://en.wikipedia.org/wiki/LaToya_London
Latrell Sprewell	http://en.wikipedia.org/wiki/Latrell_Sprewell
Laura Aikman	http://en.wikipedia.org/wiki/Laura_Aikman
Laura Antonelli	http://en.wikipedia.org/wiki/Laura_Antonelli
Laura Baugh	http://en.wikipedia.org/wiki/Laura_Baugh
Laura Branigan	http://en.wikipedia.org/wiki/Laura_Branigan
Laura Bush	http://en.wikipedia.org/wiki/Laura_Bush
Laura Chinchilla	http://en.wikipedia.org/wiki/Laura_Chinchilla
Laura Day	http://en.wikipedia.org/wiki/Laura_Day
Laura Dern	http://en.wikipedia.org/wiki/Laura_Dern
Laura Hillenbrand	http://en.wikipedia.org/wiki/Laura_Hillenbrand
Laura Ingalls Wilder	http://en.wikipedia.org/wiki/Laura_Ingalls_Wilder
Laura Ingraham	http://en.wikipedia.org/wiki/Laura_Ingraham
Laura Innes	http://en.wikipedia.org/wiki/Laura_Innes
Laura Kightlinger	http://en.wikipedia.org/wiki/Laura_Kightlinger
Laura Leighton	http://en.wikipedia.org/wiki/Laura_Leighton
Laura Linney	http://en.wikipedia.org/wiki/Laura_Linney
Laura Miller	http://en.wikipedia.org/wiki/Laura_Miller
Laura Nyro	http://en.wikipedia.org/wiki/Laura_Nyro
Laura Prepon	http://en.wikipedia.org/wiki/Laura_Prepon
Laura Richardson	http://en.wikipedia.org/wiki/Laura_Richardson
Laura Riding	http://en.wikipedia.org/wiki/Laura_Riding
Laura San Giacomo	http://en.wikipedia.org/wiki/Laura_San_Giacomo
Laura Sandys	http://en.wikipedia.org/wiki/Laura_Sandys
Laura Schlessinger	http://en.wikipedia.org/wiki/Laura_Schlessinger
Laura Z. Hobson	http://en.wikipedia.org/wiki/Laura_Z._Hobson
Laurance Rockefeller	http://en.wikipedia.org/wiki/Laurance_Rockefeller
Laurel Holloman	http://en.wikipedia.org/wiki/Laurel_Holloman
Laurell K. Hamilton	http://en.wikipedia.org/wiki/Laurell_K._Hamilton
Lauren Ambrose	http://en.wikipedia.org/wiki/Lauren_Ambrose
Lauren Anderson	http://en.wikipedia.org/wiki/Lauren_Anderson
Lauren Bacall	http://en.wikipedia.org/wiki/Lauren_Bacall
Lauren Bush	http://en.wikipedia.org/wiki/Lauren_Bush
Lauren Collins	http://en.wikipedia.org/wiki/Lauren_Collins
Lauren Graham	http://en.wikipedia.org/wiki/Lauren_Graham
Lauren Holly	http://en.wikipedia.org/wiki/Lauren_Holly
Lauren Hutton	http://en.wikipedia.org/wiki/Lauren_Hutton
Lauren Lane	http://en.wikipedia.org/wiki/Lauren_Lane
Lauren Tewes	http://en.wikipedia.org/wiki/Lauren_Tewes
Laurence Fishburne	http://en.wikipedia.org/wiki/Laurence_Fishburne
Laurence H. Meyer	http://en.wikipedia.org/wiki/Laurence_Meyer
Laurence Harvey	http://en.wikipedia.org/wiki/Laurence_Harvey
Laurence J. Peter	http://en.wikipedia.org/wiki/Laurence_J._Peter
Laurence Oliphant	http://en.wikipedia.org/wiki/Laurence_Oliphant_%28author%29
Laurence Olivier	http://en.wikipedia.org/wiki/Laurence_Olivier
Laurence Robertson	http://en.wikipedia.org/wiki/Laurence_Robertson
Laurence Sterne	http://en.wikipedia.org/wiki/Laurence_Sterne
Laurence Tisch	http://en.wikipedia.org/wiki/Laurence_Tisch
Laurence Tribe	http://en.wikipedia.org/wiki/Laurence_Tribe
Laurens Hammond	http://en.wikipedia.org/wiki/Laurens_Hammond
Laurens van der Post	http://en.wikipedia.org/wiki/Laurens_van_der_Post
Laurent Gbagbo	http://en.wikipedia.org/wiki/Laurent_Gbagbo
Lauri Ylönen	http://en.wikipedia.org/wiki/Lauri_Yl%C3%B6nen
Laurie Anderson	http://en.wikipedia.org/wiki/Laurie_Anderson
Laurie Dhue	http://en.wikipedia.org/wiki/Laurie_Dhue
Laurie Metcalf	http://en.wikipedia.org/wiki/Laurie_Metcalf
Laurie Morgan	http://en.wikipedia.org/wiki/Laurie_Morgan
Lauryn Hill	http://en.wikipedia.org/wiki/Lauryn_Hill
LaWanda Page	http://en.wikipedia.org/wiki/LaWanda_Page
Lawrence Alma-Tadema	http://en.wikipedia.org/wiki/Lawrence_Alma-Tadema
Lawrence Bragg	http://en.wikipedia.org/wiki/Lawrence_Bragg
Lawrence Coughlin	http://en.wikipedia.org/wiki/Lawrence_Coughlin
Lawrence Durrell	http://en.wikipedia.org/wiki/Lawrence_Durrell
Lawrence E. Walsh	http://en.wikipedia.org/wiki/Lawrence_E._Walsh
Lawrence Eagleburger	http://en.wikipedia.org/wiki/Lawrence_Eagleburger
Lawrence F. Probst III 	http://en.wikipedia.org/wiki/Larry_Probst
Lawrence Ferlinghetti	http://en.wikipedia.org/wiki/Lawrence_Ferlinghetti
Lawrence Gonzi	http://en.wikipedia.org/wiki/Lawrence_Gonzi
Lawrence H. Summers	http://en.wikipedia.org/wiki/Lawrence_H._Summers
Lawrence J. Korb	http://en.wikipedia.org/wiki/Lawrence_Korb
Lawrence J. Smith	http://en.wikipedia.org/wiki/Lawrence_J._Smith
Lawrence K. White	http://en.wikipedia.org/wiki/Lawrence_Kermit_White
Lawrence Kasdan	http://en.wikipedia.org/wiki/Lawrence_Kasdan
Lawrence Kudlow	http://en.wikipedia.org/wiki/Lawrence_Kudlow
Lawrence Lessig	http://en.wikipedia.org/wiki/Lawrence_Lessig
Lawrence O'Donnell	http://en.wikipedia.org/wiki/Lawrence_O%27Donnell
Lawrence Phillips	http://en.wikipedia.org/wiki/Lawrence_Phillips
Lawrence Pressman	http://en.wikipedia.org/wiki/Lawrence_Pressman
Lawrence Taylor	http://en.wikipedia.org/wiki/Lawrence_Taylor
Lawrence Tierney	http://en.wikipedia.org/wiki/Lawrence_Tierney
Lawrence Welk	http://en.wikipedia.org/wiki/Lawrence_Welk
Lawton Chiles	http://en.wikipedia.org/wiki/Lawton_Chiles
Layne Staley	http://en.wikipedia.org/wiki/Layne_Staley
Lazare Carnot	http://en.wikipedia.org/wiki/Lazare_Carnot
Lazare Hoche	http://en.wikipedia.org/wiki/Lazare_Hoche
Le Corbusier	http://en.wikipedia.org/wiki/Le_Corbusier
Le Duc Tho	http://en.wikipedia.org/wiki/Le_Duc_Tho
Lea Salonga	http://en.wikipedia.org/wiki/Lea_Salonga
Lea Thompson	http://en.wikipedia.org/wiki/Lea_Thompson
Leah Remini	http://en.wikipedia.org/wiki/Leah_Remini
Leander Starr Jameson	http://en.wikipedia.org/wiki/Leander_Starr_Jameson
LeAnn Rimes	http://en.wikipedia.org/wiki/LeAnn_Rimes
Learned Hand	http://en.wikipedia.org/wiki/Learned_Hand
LeBron James	http://en.wikipedia.org/wiki/LeBron_James
Lech Kaczynski	http://en.wikipedia.org/wiki/Lech_Kaczy%C5%84ski
Lech Walesa	http://en.wikipedia.org/wiki/Lech_Walesa
Lee "Scratch" Perry	http://en.wikipedia.org/wiki/Lee_Perry
Lee Aaker	http://en.wikipedia.org/wiki/Lee_Aaker
Lee Ann Womack	http://en.wikipedia.org/wiki/Lee_Ann_Womack
Lee Atwater	http://en.wikipedia.org/wiki/Lee_Atwater
Lee De Forest	http://en.wikipedia.org/wiki/Lee_De_Forest
Lee Grant	http://en.wikipedia.org/wiki/Lee_Grant
Lee Greenwood	http://en.wikipedia.org/wiki/Lee_Greenwood
Lee H. Hamilton	http://en.wikipedia.org/wiki/Lee_H._Hamilton
Lee Hai-chan	http://en.wikipedia.org/wiki/Lee_Hai-chan
Lee Harvey Oswald	http://en.wikipedia.org/wiki/Lee_Harvey_Oswald
Lee Hazlewood	http://en.wikipedia.org/wiki/Lee_Hazlewood
Lee Horsley	http://en.wikipedia.org/wiki/Lee_Horsley
Lee Hsien Loong	http://en.wikipedia.org/wiki/Lee_Hsien_Loong
Lee Iacocca	http://en.wikipedia.org/wiki/Lee_Iacocca
Lee J. Cobb	http://en.wikipedia.org/wiki/Lee_J._Cobb
Lee Jong-Wook	http://en.wikipedia.org/wiki/Lee_Jong-wook
Lee Krasner	http://en.wikipedia.org/wiki/Lee_Krasner
Lee Kuan Yew	http://en.wikipedia.org/wiki/Lee_Kuan_Yew
Lee Majors	http://en.wikipedia.org/wiki/Lee_Majors
Lee Malvo	http://en.wikipedia.org/wiki/Lee_Malvo
Lee Marvin	http://en.wikipedia.org/wiki/Lee_Marvin
Lee Meriwether	http://en.wikipedia.org/wiki/Lee_Meriwether
Lee Myung-bak	http://en.wikipedia.org/wiki/Lee_Myung-bak
Lee Patrick	http://en.wikipedia.org/wiki/Lee_Patrick_%28actress%29
Lee R. Raymond	http://en.wikipedia.org/wiki/Lee_R._Raymond
Lee Radziwill	http://en.wikipedia.org/wiki/Lee_Radziwill
Lee Remick	http://en.wikipedia.org/wiki/Lee_Remick
Lee Ritenour	http://en.wikipedia.org/wiki/Lee_Ritenour
Lee Ryan	http://en.wikipedia.org/wiki/Lee_Ryan
Lee Scott	http://en.wikipedia.org/wiki/Lee_Scott_%28UK_politician%29
Lee Smith	http://en.wikipedia.org/wiki/Lee_Smith_%28fiction_author%29
Lee Strasberg	http://en.wikipedia.org/wiki/Lee_Strasberg
Lee Tamahori	http://en.wikipedia.org/wiki/Lee_Tamahori
Lee Tergesen	http://en.wikipedia.org/wiki/Lee_Tergesen
Lee Terry	http://en.wikipedia.org/wiki/Lee_Terry
Lee Tracy	http://en.wikipedia.org/wiki/Lee_Tracy
Lee Trevino	http://en.wikipedia.org/wiki/Lee_Trevino
Lee Van Cleef	http://en.wikipedia.org/wiki/Lee_Van_Cleef
Leelee Sobieski	http://en.wikipedia.org/wiki/Leelee_Sobieski
Leeza Gibbons	http://en.wikipedia.org/wiki/Leeza_Gibbons
Lefty Grove	http://en.wikipedia.org/wiki/Lefty_Grove
Legs Larry Smith	http://en.wikipedia.org/wiki/Larry_Smith_(musician)
Leif Erickson	http://en.wikipedia.org/wiki/Leif_Erickson
Leif Ericsson	http://en.wikipedia.org/wiki/Leif_Ericson
Leif Garrett	http://en.wikipedia.org/wiki/Leif_Garrett
Leigh Hunt	http://en.wikipedia.org/wiki/Leigh_Hunt
Leigh McCloskey	http://en.wikipedia.org/wiki/Leigh_McCloskey
Leigh Taylor-Young	http://en.wikipedia.org/wiki/Leigh_Taylor-Young
Leighton Meesters	http://en.wikipedia.org/wiki/Leighton_Meester
Leisha Hailey	http://en.wikipedia.org/wiki/Leisha_Hailey
Lela Rochon	http://en.wikipedia.org/wiki/Lela_Rochon
Leland Chapman	http://en.wikipedia.org/wiki/Leland_Chapman
Leland Stanford	http://en.wikipedia.org/wiki/Leland_Stanford
Leland Yee	http://en.wikipedia.org/wiki/Leland_Yee
Lemony Snicket	http://en.wikipedia.org/wiki/Lemony_Snicket
Len Dawson	http://en.wikipedia.org/wiki/Len_Dawson
Len Deighton	http://en.wikipedia.org/wiki/Len_Deighton
Lena Horne	http://en.wikipedia.org/wiki/Lena_Horne
Lena Katina	http://en.wikipedia.org/wiki/Lena_Katina
Lena Olin	http://en.wikipedia.org/wiki/Lena_Olin
Leni Riefenstahl	http://en.wikipedia.org/wiki/Leni_Riefenstahl
Lennart Meri	http://en.wikipedia.org/wiki/Lennart_Meri
Lennox Lewis	http://en.wikipedia.org/wiki/Lennox_Lewis
Lenny Bruce	http://en.wikipedia.org/wiki/Lenny_Bruce
Lenny Henry	http://en.wikipedia.org/wiki/Lenny_Henry
Lenny Kravitz	http://en.wikipedia.org/wiki/Lenny_Kravitz
Lenny Wilkens	http://en.wikipedia.org/wiki/Lenny_Wilkens
Leo Baekeland	http://en.wikipedia.org/wiki/Leo_Baekeland
Leo Burnett	http://en.wikipedia.org/wiki/Leo_Burnett
Leo Buscaglia	http://en.wikipedia.org/wiki/Leo_Buscaglia
L�o Delibes	http://en.wikipedia.org/wiki/L%e9o_Delibes
Leo Durocher	http://en.wikipedia.org/wiki/Leo_Durocher
Leo Esaki	http://en.wikipedia.org/wiki/Leo_Esaki
Leo Fender	http://en.wikipedia.org/wiki/Leo_Fender
Leo G. Carroll	http://en.wikipedia.org/wiki/Leo_G._Carroll
Leo Gorcey	http://en.wikipedia.org/wiki/Leo_Gorcey
Leo Kottke	http://en.wikipedia.org/wiki/Leo_Kottke
Leo Laporte	http://en.wikipedia.org/wiki/Leo_Laporte
Leo McCarey	http://en.wikipedia.org/wiki/Leo_McCarey
Leo McKern	http://en.wikipedia.org/wiki/Leo_McKern
Leo Penn	http://en.wikipedia.org/wiki/Leo_Penn
Leo Rosten	http://en.wikipedia.org/wiki/Leo_Rosten
Leo Ryan	http://en.wikipedia.org/wiki/Leo_Ryan
Leo Sayer	http://en.wikipedia.org/wiki/Leo_Sayer
Leo Strauss	http://en.wikipedia.org/wiki/Leo_Strauss
Leo Szilard	http://en.wikipedia.org/wiki/Le%C3%B3_Szil%C3%A1rd
Leo Tolstoy	http://en.wikipedia.org/wiki/Leo_Tolstoy
Leo von Caprivi	http://en.wikipedia.org/wiki/Leo_von_Caprivi
Leo XIII	http://en.wikipedia.org/wiki/Leo_XIII
Leon Ames	http://en.wikipedia.org/wiki/Leon_Ames_%28actor%29
Leon Askin	http://en.wikipedia.org/wiki/Leon_Askin
Leon Battista Alberti	http://en.wikipedia.org/wiki/Leon_Battista_Alberti
L�on Bourgeois	http://en.wikipedia.org/wiki/L%e9on_Bourgeois
Leon Czolgosz	http://en.wikipedia.org/wiki/Leon_Czolgosz
Leon Edel	http://en.wikipedia.org/wiki/Leon_Edel
L�on Foucault	http://en.wikipedia.org/wiki/L%e9on_Foucault
L�on Gambetta	http://en.wikipedia.org/wiki/L%e9on_Gambetta
Leon Jaworski	http://en.wikipedia.org/wiki/Leon_Jaworski
Leon Jouhaux	http://en.wikipedia.org/wiki/L%C3%A9on_Jouhaux
Leon Klinghoffer	http://en.wikipedia.org/wiki/Leon_Klinghoffer
Leon M. Lederman	http://en.wikipedia.org/wiki/Leon_M._Lederman
Leon N. Cooper	http://en.wikipedia.org/wiki/Leon_N._Cooper
Leon of Modena	http://en.wikipedia.org/wiki/Leon_of_Modena
Leon Panetta	http://en.wikipedia.org/wiki/Leon_Panetta
Leon Redbone	http://en.wikipedia.org/wiki/Leon_Redbone
Leon Russell	http://en.wikipedia.org/wiki/Leon_Russell
Leon Spinks	http://en.wikipedia.org/wiki/Leon_Spinks
Leon Trotsky	http://en.wikipedia.org/wiki/Leon_Trotsky
Leon Uris	http://en.wikipedia.org/wiki/Leon_Uris
L�on Walras	http://en.wikipedia.org/wiki/L%e9on_Walras
Leon Wieseltier	http://en.wikipedia.org/wiki/Leon_Wieseltier
Leona Helmsley	http://en.wikipedia.org/wiki/Leona_Helmsley
Leonard Baskin	http://en.wikipedia.org/wiki/Leonard_Baskin
Leonard Bernstein	http://en.wikipedia.org/wiki/Leonard_Bernstein
Leonard Boswell	http://en.wikipedia.org/wiki/Leonard_Boswell
Leonard Carmichael	http://en.wikipedia.org/wiki/Leonard_Carmichael
Leonard Cohen	http://en.wikipedia.org/wiki/Leonard_Cohen
Leonard Horner	http://en.wikipedia.org/wiki/Leonard_Horner
Leonard Lance	http://en.wikipedia.org/wiki/Leonard_Lance
Leonard Little	http://en.wikipedia.org/wiki/Leonard_Little
Leonard Maltin	http://en.wikipedia.org/wiki/Leonard_Maltin
Leonard Nimoy	http://en.wikipedia.org/wiki/Leonard_Nimoy
Leonard Peikoff	http://en.wikipedia.org/wiki/Leonard_Peikoff
Leonard Peltier	http://en.wikipedia.org/wiki/Leonard_Peltier
Leonard Rossiter	http://en.wikipedia.org/wiki/Leonard_Rossiter
Leonard Stern	http://en.wikipedia.org/wiki/Leonard_N._Stern
Leonard Whiting	http://en.wikipedia.org/wiki/Leonard_Whiting
Leonard Woodcock	http://en.wikipedia.org/wiki/Leonard_Woodcock
Leonard Woolf	http://en.wikipedia.org/wiki/Leonard_Woolf
Leonardo Da Vinci	http://en.wikipedia.org/wiki/Leonardo_da_Vinci
Leonardo DiCaprio	http://en.wikipedia.org/wiki/Leonardo_DiCaprio
Leonardo Fibonacci	http://en.wikipedia.org/wiki/Leonardo_Fibonacci
Leonel Fern�ndez	http://en.wikipedia.org/wiki/Leonel_Fern%C3%A1ndez
Leonhard Euler	http://en.wikipedia.org/wiki/Leonhard_Euler
Leonid Brezhnev	http://en.wikipedia.org/wiki/Leonid_Brezhnev
Leonid Kuchma	http://en.wikipedia.org/wiki/Leonid_Kuchma
Leonidas Polk	http://en.wikipedia.org/wiki/Leonidas_Polk
L�onie Adams	http://en.wikipedia.org/wiki/L%e9onie_Adams
Leonor Fini	http://en.wikipedia.org/wiki/Leonor_Fini
Leontyne Price	http://en.wikipedia.org/wiki/Leontyne_Price
Leopold I	http://en.wikipedia.org/wiki/Leopold_I_of_Belgium
Leopold II	http://en.wikipedia.org/wiki/Leopold_II_of_Belgium
Leopold III	http://en.wikipedia.org/wiki/Leopold_III_of_Belgium
Leopold Ruzicka	http://en.wikipedia.org/wiki/Leopold_Ru%C5%BEi%C4%8Dka
L�opold Senghor	http://en.wikipedia.org/wiki/L%e9opold_Senghor
Leopold von Ranke	http://en.wikipedia.org/wiki/Leopold_von_Ranke
Leopoldo Galtieri	http://en.wikipedia.org/wiki/Leopoldo_Galtieri
Leo� Jan�cek	http://en.wikipedia.org/wiki/Leo%C5%A1_Jan%C3%A1%C4%8Dek
Leroy Anderson	http://en.wikipedia.org/wiki/Leroy_Anderson
Leroy Burrell	http://en.wikipedia.org/wiki/Leroy_Burrell
Leroy Grumman	http://en.wikipedia.org/wiki/Leroy_Grumman
Les Aspin	http://en.wikipedia.org/wiki/Les_Aspin
Les AuCoin	http://en.wikipedia.org/wiki/Les_AuCoin
Les Baxter	http://en.wikipedia.org/wiki/Les_Baxter
Les Brown	http://en.wikipedia.org/wiki/Les_Brown_%28bandleader%29
Les Claypool	http://en.wikipedia.org/wiki/Les_Claypool
Les Moonves	http://en.wikipedia.org/wiki/Les_Moonves
Les Paul	http://en.wikipedia.org/wiki/Les_Paul
Les Tremayne	http://en.wikipedia.org/wiki/Les_Tremayne
Lesley Ann Warren	http://en.wikipedia.org/wiki/Lesley_Ann_Warren
Lesley Boone	http://en.wikipedia.org/wiki/Lesley_Boone
Lesley Gore	http://en.wikipedia.org/wiki/Lesley_Gore
Lesley Stahl	http://en.wikipedia.org/wiki/Lesley_Stahl
Lesley-Anne Down	http://en.wikipedia.org/wiki/Lesley-Anne_Down
Leslie A. Fiedler	http://en.wikipedia.org/wiki/Leslie_A._Fiedler
Leslie A. White	http://en.wikipedia.org/wiki/Leslie_A._White
Leslie Banks	http://en.wikipedia.org/wiki/Leslie_Banks
Leslie Caron	http://en.wikipedia.org/wiki/Leslie_Caron
Leslie Charteris	http://en.wikipedia.org/wiki/Leslie_Charteris
Leslie Easterbrook	http://en.wikipedia.org/wiki/Leslie_Easterbrook
Leslie H. Gelb	http://en.wikipedia.org/wiki/Leslie_H._Gelb
Leslie Howard	http://en.wikipedia.org/wiki/Leslie_Howard_%28actor%29
Leslie Jordan	http://en.wikipedia.org/wiki/Leslie_Jordan
Leslie Nielsen	http://en.wikipedia.org/wiki/Leslie_Nielsen
Leslie R. Groves	http://en.wikipedia.org/wiki/Leslie_R._Groves
Leslie Uggams	http://en.wikipedia.org/wiki/Leslie_Uggams
Lester Bangs	http://en.wikipedia.org/wiki/Lester_Bangs
Lester Bowie	http://en.wikipedia.org/wiki/Lester_Bowie
Lester Bowles Pearson	http://en.wikipedia.org/wiki/Lester_Bowles_Pearson
Lester Crawford	http://en.wikipedia.org/wiki/Lester_Crawford
Lester del Rey	http://en.wikipedia.org/wiki/Lester_del_Rey
Lester Maddox	http://en.wikipedia.org/wiki/Lester_Maddox
Lester Thurow	http://en.wikipedia.org/wiki/Lester_Thurow
Lester Young	http://en.wikipedia.org/wiki/Lester_Young
Letsie III	http://en.wikipedia.org/wiki/Letsie_III_of_Lesotho
Lev Landau	http://en.wikipedia.org/wiki/Lev_Landau
Lev Yashin	http://en.wikipedia.org/wiki/Lev_Yashin
LeVar Burton	http://en.wikipedia.org/wiki/LeVar_Burton
Leverett Saltonstall	http://en.wikipedia.org/wiki/Leverett_Saltonstall
Levi Eshkol	http://en.wikipedia.org/wiki/Levi_Eshkol
Levi P. Morton	http://en.wikipedia.org/wiki/Levi_P._Morton
Levon Helm	http://en.wikipedia.org/wiki/Levon_Helm
Levy Mwanawasa	http://en.wikipedia.org/wiki/Levy_Mwanawasa
Lew Ayres	http://en.wikipedia.org/wiki/Lew_Ayres
Lew Wallace	http://en.wikipedia.org/wiki/Lew_Wallace
Lew Wasserman	http://en.wikipedia.org/wiki/Lew_Wasserman
Lewis B. Hershey	http://en.wikipedia.org/wiki/Lewis_B._Hershey
Lewis Black	http://en.wikipedia.org/wiki/Lewis_Black
Lewis Carroll	http://en.wikipedia.org/wiki/Lewis_Carroll
Lewis Cass	http://en.wikipedia.org/wiki/Lewis_Cass
Lewis F. Powell, Jr.	http://en.wikipedia.org/wiki/Lewis_F._Powell,_Jr.
Lewis Gilbert	http://en.wikipedia.org/wiki/Lewis_Gilbert
Lewis Henry Morgan	http://en.wikipedia.org/wiki/Lewis_Henry_Morgan
Lewis Libby	http://en.wikipedia.org/wiki/Lewis_Libby
Lewis Milestone	http://en.wikipedia.org/wiki/Lewis_Milestone
Lewis Mumford	http://en.wikipedia.org/wiki/Lewis_Mumford
Lewis Seiler	http://en.wikipedia.org/wiki/Lewis_Seiler
Lewis Stone	http://en.wikipedia.org/wiki/Lewis_Stone
Lewis Teague	http://en.wikipedia.org/wiki/Lewis_Teague
Lex Barker	http://en.wikipedia.org/wiki/Lex_Barker
Lexa Doig	http://en.wikipedia.org/wiki/Lexa_Doig
Li Gong	http://en.wikipedia.org/wiki/Gong_Li
Liam Aiken	http://en.wikipedia.org/wiki/Liam_Aiken
Liam Byrne	http://en.wikipedia.org/wiki/Liam_Byrne
Liam Fox	http://en.wikipedia.org/wiki/Liam_Fox
Liam Gallagher	http://en.wikipedia.org/wiki/Liam_Gallagher
Liam Howlett	http://en.wikipedia.org/wiki/Liam_Howlett
Liam Neeson	http://en.wikipedia.org/wiki/Liam_Neeson
Liam O'Flaherty	http://en.wikipedia.org/wiki/Liam_O%27Flaherty
Lieutenant-General Soe Win	http://en.wikipedia.org/wiki/Soe_Win
Liev Schreiber	http://en.wikipedia.org/wiki/Liev_Schreiber
Lil' Fizz	http://en.wikipedia.org/wiki/Lil%27_Fizz
Lil' Flip	http://en.wikipedia.org/wiki/Lil%27_Flip
Lil' Jon	http://en.wikipedia.org/wiki/Lil%27_Jon
Lil' Kim	http://en.wikipedia.org/wiki/Lil%27_Kim
Lil' Mo	http://en.wikipedia.org/wiki/Lil%27_Mo
Lil' Rob	http://en.wikipedia.org/wiki/Lil_Rob
Lil' Romeo	http://en.wikipedia.org/wiki/Lil%27_Romeo
Lil' Scrappy	http://en.wikipedia.org/wiki/Lil_Scrappy
Lil' Wayne	http://en.wikipedia.org/wiki/Lil_Wayne
Lila Kedrova	http://en.wikipedia.org/wiki/Lila_Kedrova
Lila Wallace	http://en.wikipedia.org/wiki/Lila_Wallace
Lili Damita	http://en.wikipedia.org/wiki/Lili_Damita
Lili Taylor	http://en.wikipedia.org/wiki/Lili_Taylor
Lilian Greenwood	http://en.wikipedia.org/wiki/Lilian_Greenwood
Liliana Abud	http://en.wikipedia.org/wiki/Liliana_Abud
Liliane Bettencourt	http://en.wikipedia.org/wiki/Liliane_Bettencourt
Lilli Palmer	http://en.wikipedia.org/wiki/Lilli_Palmer
Lillian Gish	http://en.wikipedia.org/wiki/Lillian_Gish
Lillian Hellman	http://en.wikipedia.org/wiki/Lillian_Hellman
Lillian Roth	http://en.wikipedia.org/wiki/Lillian_Roth
Lillie Hitchcock Coit	http://en.wikipedia.org/wiki/Lillie_Hitchcock_Coit
Lillo Brancato	http://en.wikipedia.org/wiki/Lillo_Brancato,_Jr.
Lily Tomlin	http://en.wikipedia.org/wiki/Lily_Tomlin
Lilyan Tashman	http://en.wikipedia.org/wiki/Lilyan_Tashman
Lina Wertmüller	http://en.wikipedia.org/wiki/Lina_Wertm%C3%BCller
Lincoln Chafee	http://en.wikipedia.org/wiki/Lincoln_Chafee
Lincoln Davis	http://en.wikipedia.org/wiki/Lincoln_Davis
Lincoln Diaz-Balart	http://en.wikipedia.org/wiki/Lincoln_Diaz-Balart
Lincoln Kirstein	http://en.wikipedia.org/wiki/Lincoln_Kirstein
Lincoln Steffens	http://en.wikipedia.org/wiki/Lincoln_Steffens
Linda Blair	http://en.wikipedia.org/wiki/Linda_Blair
Linda Cardellini	http://en.wikipedia.org/wiki/Linda_Cardellini
Linda Chavez	http://en.wikipedia.org/wiki/Linda_Chavez
Linda Darnell	http://en.wikipedia.org/wiki/Linda_Darnell
Linda Ellerbee	http://en.wikipedia.org/wiki/Linda_Ellerbee
Linda Evangelista	http://en.wikipedia.org/wiki/Linda_Evangelista
Linda Evans	http://en.wikipedia.org/wiki/Linda_Evans
Linda Fiorentino	http://en.wikipedia.org/wiki/Linda_Fiorentino
Linda Gray	http://en.wikipedia.org/wiki/Linda_Gray
Linda Hamilton	http://en.wikipedia.org/wiki/Linda_Hamilton
Linda Hunt	http://en.wikipedia.org/wiki/Linda_Hunt
Linda Kelsey	http://en.wikipedia.org/wiki/Linda_Kelsey
Linda Kozlowski	http://en.wikipedia.org/wiki/Linda_Kozlowski
Linda Lavin	http://en.wikipedia.org/wiki/Linda_Lavin
Linda Lingle	http://en.wikipedia.org/wiki/Linda_Lingle
Linda McCartney	http://en.wikipedia.org/wiki/Linda_McCartney
Linda Perry	http://en.wikipedia.org/wiki/Linda_Perry
Linda Purl	http://en.wikipedia.org/wiki/Linda_Purl
Linda Riordan	http://en.wikipedia.org/wiki/Linda_Riordan
Linda Ronstadt	http://en.wikipedia.org/wiki/Linda_Ronstadt
Linda S�nchez	http://en.wikipedia.org/wiki/Linda_S%C3%A1nchez
Linda Tripp	http://en.wikipedia.org/wiki/Linda_Tripp
Linda Vester	http://en.wikipedia.org/wiki/Linda_Vester
Lindsay Anderson	http://en.wikipedia.org/wiki/Lindsay_Anderson
Lindsay Crosby	http://en.wikipedia.org/wiki/Lindsay_Crosby
Lindsay Crouse	http://en.wikipedia.org/wiki/Lindsay_Crouse
Lindsay Hoyle	http://en.wikipedia.org/wiki/Lindsay_Hoyle
Lindsay Kemp	http://en.wikipedia.org/wiki/Lindsay_Kemp
Lindsay Lohan	http://en.wikipedia.org/wiki/Lindsay_Lohan
Lindsay Owen-Jones	http://en.wikipedia.org/wiki/Lindsay_Owen-Jones
Lindsay Price	http://en.wikipedia.org/wiki/Lindsay_Price
Lindsay Roy	http://en.wikipedia.org/wiki/Lindsay_Roy
Lindsay Thomas	http://en.wikipedia.org/wiki/Lindsay_Thomas_%28politician%29
Lindsay Wagner	http://en.wikipedia.org/wiki/Lindsay_Wagner
Lindsey Buckingham	http://en.wikipedia.org/wiki/Lindsey_Buckingham
Lindsey Graham	http://en.wikipedia.org/wiki/Lindsey_Graham
Lindy Boggs	http://en.wikipedia.org/wiki/Lindy_Boggs
Link Wray	http://en.wikipedia.org/wiki/Link_Wray
Linus Pauling	http://en.wikipedia.org/wiki/Linus_Pauling
Linus Torvalds	http://en.wikipedia.org/wiki/Linus_Torvalds
Lionel Atwill	http://en.wikipedia.org/wiki/Lionel_Atwill
Lionel Barrymore	http://en.wikipedia.org/wiki/Lionel_Barrymore
Lionel Hampton	http://en.wikipedia.org/wiki/Lionel_Hampton
Lionel Jeffries	http://en.wikipedia.org/wiki/Lionel_Jeffries
Lionel Jospin	http://en.wikipedia.org/wiki/Lionel_Jospin
Lionel Richie	http://en.wikipedia.org/wiki/Lionel_Richie
Lionel Stander	http://en.wikipedia.org/wiki/Lionel_Stander
Lionel Tate	http://en.wikipedia.org/wiki/Lionel_Tate
Lionel Tiger	http://en.wikipedia.org/wiki/Lionel_Tiger
Lionel Trilling	http://en.wikipedia.org/wiki/Lionel_Trilling
Lisa "Left Eye" Lopes	http://en.wikipedia.org/wiki/Lisa_%22Left_Eye%22_Lopes
Lisa Blount	http://en.wikipedia.org/wiki/Lisa_Blount
Lisa Bonet	http://en.wikipedia.org/wiki/Lisa_Bonet
Lisa Boyle	http://en.wikipedia.org/wiki/Lisa_Boyle
Lisa Carver	http://en.wikipedia.org/wiki/Lisa_Carver
Lisa Daniels	http://en.wikipedia.org/wiki/Lisa_Daniels_%28TV_presenter%29
Lisa Edelstein	http://en.wikipedia.org/wiki/Lisa_Edelstein
Lisa Hartman	http://en.wikipedia.org/wiki/Lisa_Hartman
Lisa Kudrow	http://en.wikipedia.org/wiki/Lisa_Kudrow
Lisa Leslie	http://en.wikipedia.org/wiki/Lisa_Leslie
Lisa Loeb	http://en.wikipedia.org/wiki/Lisa_Loeb
Lisa Loring	http://en.wikipedia.org/wiki/Lisa_Loring
Lisa Marie Presley	http://en.wikipedia.org/wiki/Lisa_Marie_Presley
Lisa Murkowski	http://en.wikipedia.org/wiki/Lisa_Murkowski
Lisa Nandy	http://en.wikipedia.org/wiki/Lisa_Nandy
Lisa Nicole Carson	http://en.wikipedia.org/wiki/Lisa_Nicole_Carson
Lisa Raye	http://en.wikipedia.org/wiki/Lisa_Raye
Lisa Rinna	http://en.wikipedia.org/wiki/Lisa_Rinna
Lisa Whelchel	http://en.wikipedia.org/wiki/Lisa_Whelchel
Lise Meitner	http://en.wikipedia.org/wiki/Lise_Meitner
Lisel Mueller	http://en.wikipedia.org/wiki/Lisel_Mueller
Lita Ford	http://en.wikipedia.org/wiki/Lita_Ford
Little Eva	http://en.wikipedia.org/wiki/Little_Eva
Little Jimmy Dickens	http://en.wikipedia.org/wiki/Little_Jimmy_Dickens
Little Milton	http://en.wikipedia.org/wiki/Little_Milton
Little Richard	http://en.wikipedia.org/wiki/Little_Richard
Little Willie John	http://en.wikipedia.org/wiki/Little_Willie_John
Liv Tyler	http://en.wikipedia.org/wiki/Liv_Tyler
Liv Ullmann	http://en.wikipedia.org/wiki/Liv_Ullmann
Livia Drusilla	http://en.wikipedia.org/wiki/Livia_Drusilla
Liz Claiborne	http://en.wikipedia.org/wiki/Liz_Claiborne_%28fashion_designer%29
Liz Phair	http://en.wikipedia.org/wiki/Liz_Phair
Liza Minnelli	http://en.wikipedia.org/wiki/Liza_Minnelli
Lizabeth Scott	http://en.wikipedia.org/wiki/Lizabeth_Scott
Lizette Woodworth Reese	http://en.wikipedia.org/wiki/Lizette_Woodworth_Reese
Lizzie Grubman	http://en.wikipedia.org/wiki/Lizzie_Grubman
Ljubco Georgievski	http://en.wikipedia.org/wiki/Ljub%C4%8Do_Georgievski
LL Cool J	http://en.wikipedia.org/wiki/LL_Cool_J
Lleyton Hewitt	http://en.wikipedia.org/wiki/Lleyton_Hewitt
Lloyd Alexander	http://en.wikipedia.org/wiki/Lloyd_Alexander
Lloyd Bacon	http://en.wikipedia.org/wiki/Lloyd_Bacon
Lloyd Banks	http://en.wikipedia.org/wiki/Lloyd_Banks
Lloyd Bentsen, Jr.	http://en.wikipedia.org/wiki/Lloyd_Bentsen
Lloyd Blankfein	http://en.wikipedia.org/wiki/Lloyd_Blankfein
Lloyd Bochner	http://en.wikipedia.org/wiki/Lloyd_Bochner
Lloyd Bridges	http://en.wikipedia.org/wiki/Lloyd_Bridges
Lloyd Bucher	http://en.wikipedia.org/wiki/Lloyd_Bucher
Lloyd Doggett	http://en.wikipedia.org/wiki/Lloyd_Doggett
Lloyd Gough	http://en.wikipedia.org/wiki/Lloyd_Gough
Lloyd Kaufman	http://en.wikipedia.org/wiki/Lloyd_Kaufman
Lloyd Meeds	http://en.wikipedia.org/wiki/Lloyd_Meeds
Lois Capps	http://en.wikipedia.org/wiki/Lois_Capps
Lois Duncan	http://en.wikipedia.org/wiki/Lois_Duncan
Lois McMaster Bujold	http://en.wikipedia.org/wiki/Lois_McMaster_Bujold
Lol Coxhill	http://en.wikipedia.org/wiki/Lol_Coxhill
Lola Albright	http://en.wikipedia.org/wiki/Lola_Albright
Lola Montez	http://en.wikipedia.org/wiki/Lola_Montez
Lolita Davidovich	http://en.wikipedia.org/wiki/Lolita_Davidovich
Lon Chaney	http://en.wikipedia.org/wiki/Lon_Chaney,_Sr.
Lon Chaney, Jr.	http://en.wikipedia.org/wiki/Lon_Chaney,_Jr.
Lon Horiuchi	http://en.wikipedia.org/wiki/Lon_Horiuchi
Long John Baldry	http://en.wikipedia.org/wiki/Long_John_Baldry
Loni Anderson	http://en.wikipedia.org/wiki/Loni_Anderson
Lonnie Johnson	http://en.wikipedia.org/wiki/Lonnie_Johnson_%28inventor%29
Lope de Vega	http://en.wikipedia.org/wiki/Lope_de_Vega
Lord Acton	http://en.wikipedia.org/wiki/Lord_Acton
Lord Beaverbrook	http://en.wikipedia.org/wiki/Lord_Beaverbrook
Lord British	http://en.wikipedia.org/wiki/Richard_Garriott
Lord Byron	http://en.wikipedia.org/wiki/Lord_Byron
Lord Darnley	http://en.wikipedia.org/wiki/Lord_Darnley
Lord Haw-Haw	http://en.wikipedia.org/wiki/William_Joyce
Lord Kelvin	http://en.wikipedia.org/wiki/Lord_Kelvin
Lord Mountbatten	http://en.wikipedia.org/wiki/Lord_Mountbatten
Lord Nelson	http://en.wikipedia.org/wiki/Lord_Nelson
Lord Palmerston	http://en.wikipedia.org/wiki/Lord_Palmerston
Lord Randolph Churchill	http://en.wikipedia.org/wiki/Lord_Randolph_Churchill
Lord Rayleigh	http://en.wikipedia.org/wiki/Lord_Rayleigh
Lord Robertson	http://en.wikipedia.org/wiki/George_Robertson,_Baron_Robertson_of_Port_Ellen
Lorely Burt	http://en.wikipedia.org/wiki/Lorely_Burt
Loren Eiseley	http://en.wikipedia.org/wiki/Loren_Eiseley
Lorenz Hart	http://en.wikipedia.org/wiki/Lorenz_Hart
Lorenzo Bellini	http://en.wikipedia.org/wiki/Lorenzo_Bellini
Lorenzo de Medici	http://en.wikipedia.org/wiki/Lorenzo_de%27_Medici
Lorenzo di Credi	http://en.wikipedia.org/wiki/Lorenzo_di_Credi
Lorenzo Ghiberti	http://en.wikipedia.org/wiki/Lorenzo_Ghiberti
Lorenzo Lamas	http://en.wikipedia.org/wiki/Lorenzo_Lamas
Lorenzo Valla	http://en.wikipedia.org/wiki/Lorenzo_Valla
Loretta Devine	http://en.wikipedia.org/wiki/Loretta_Devine
Loretta Lynn	http://en.wikipedia.org/wiki/Loretta_Lynn
Loretta Sanchez	http://en.wikipedia.org/wiki/Loretta_Sanchez
Loretta Swit	http://en.wikipedia.org/wiki/Loretta_Swit
Loretta Young	http://en.wikipedia.org/wiki/Loretta_Young
Lori Loughlin	http://en.wikipedia.org/wiki/Lori_Loughlin
Lori Petty	http://en.wikipedia.org/wiki/Lori_Petty
Lori Singer	http://en.wikipedia.org/wiki/Lori_Singer
Lorna Luft	http://en.wikipedia.org/wiki/Lorna_Luft
Lorne Greene	http://en.wikipedia.org/wiki/Lorne_Greene
Lorne Michaels	http://en.wikipedia.org/wiki/Lorne_Michaels
Lorraine Bracco	http://en.wikipedia.org/wiki/Lorraine_Bracco
Lorraine Fullbrook	http://en.wikipedia.org/wiki/Lorraine_Fullbrook
Lorraine Hansberry	http://en.wikipedia.org/wiki/Lorraine_Hansberry
Lorraine Hunt	http://en.wikipedia.org/wiki/Lorraine_Hunt
Lothar Matth�us	http://en.wikipedia.org/wiki/Lothar_Matth%C3%A4us
Lou Adler	http://en.wikipedia.org/wiki/Lou_Adler
Lou Brock	http://en.wikipedia.org/wiki/Lou_Brock
Lou Costello	http://en.wikipedia.org/wiki/Lou_Costello
Lou Diamond Phillips	http://en.wikipedia.org/wiki/Lou_Diamond_Phillips
Lou Dobbs	http://en.wikipedia.org/wiki/Lou_Dobbs
Lou Ferrigno	http://en.wikipedia.org/wiki/Lou_Ferrigno
Lou Gehrig	http://en.wikipedia.org/wiki/Lou_Gehrig
Lou Gossett, Jr.	http://en.wikipedia.org/wiki/Lou_Gossett
Lou Gramm	http://en.wikipedia.org/wiki/Lou_Gramm
Lou Montulli	http://en.wikipedia.org/wiki/Lou_Montulli
Lou Rawls	http://en.wikipedia.org/wiki/Lou_Rawls
Lou Reed	http://en.wikipedia.org/wiki/Lou_Reed
Lou Sheldon	http://en.wikipedia.org/wiki/Lou_Sheldon
Loudon Wainwright III	http://en.wikipedia.org/wiki/Loudon_Wainwright_III
Louie Anderson	http://en.wikipedia.org/wiki/Louie_Anderson
Louie Gohmert	http://en.wikipedia.org/wiki/Louie_Gohmert
Louis A. Johnson	http://en.wikipedia.org/wiki/Louis_A._Johnson
Louis Adamic	http://en.wikipedia.org/wiki/Louis_Adamic
Louis Agassiz	http://en.wikipedia.org/wiki/Louis_Agassiz
Louis Alexandre Berthier	http://en.wikipedia.org/wiki/Louis_Alexandre_Berthier
Louis Aragon	http://en.wikipedia.org/wiki/Louis_Aragon
Louis Armstrong	http://en.wikipedia.org/wiki/Louis_Armstrong
Louis Auchincloss	http://en.wikipedia.org/wiki/Louis_Auchincloss
Louis B. Mayer	http://en.wikipedia.org/wiki/Louis_B_Mayer
Louis Braille	http://en.wikipedia.org/wiki/Louis_Braille
Louis Calhern	http://en.wikipedia.org/wiki/Louis_Calhern
Louis Christophe Fran�ois Hachette	http://en.wikipedia.org/wiki/Louis_Christophe_Fran%C3%A7ois_Hachette
Louis Comfort Tiffany	http://en.wikipedia.org/wiki/Louis_Comfort_Tiffany
Louis D. Brandeis	http://en.wikipedia.org/wiki/Louis_D._Brandeis
Louis Daguerre	http://en.wikipedia.org/wiki/Louis_Daguerre
Louis de Broglie	http://en.wikipedia.org/wiki/Louis_de_Broglie
Louis de Fun�s	http://en.wikipedia.org/wiki/Louis_de_Fun%C3%A8s
Louis Durey	http://en.wikipedia.org/wiki/Louis_Durey
Louis Farrakhan	http://en.wikipedia.org/wiki/Louis_Farrakhan
Louis Freeh	http://en.wikipedia.org/wiki/Louis_Freeh
Louis Gabriel Suchet	http://en.wikipedia.org/wiki/Louis_Gabriel_Suchet
Louis Gossett Jr.	http://en.wikipedia.org/wiki/Louis_Gossett,_Jr.
Louis Harris	http://en.wikipedia.org/wiki/Louis_Harris
Louis Hayward	http://en.wikipedia.org/wiki/Louis_Hayward
Louis Hippolyte LaFontaine	http://en.wikipedia.org/wiki/Louis-Hippolyte_Lafontaine
Louis III	http://en.wikipedia.org/wiki/Louis_III_of_France
Louis IV	http://en.wikipedia.org/wiki/Louis_IV_of_France
Louis IX	http://en.wikipedia.org/wiki/Louis_IX_of_France
Louis Jourdan	http://en.wikipedia.org/wiki/Louis_Jourdan
Louis Kahn	http://en.wikipedia.org/wiki/Louis_Kahn
Louis King	http://en.wikipedia.org/wiki/Louis_King
Louis L'Amour	http://en.wikipedia.org/wiki/Louis_L%27Amour
Louis Le Vau	http://en.wikipedia.org/wiki/Louis_Le_Vau
Louis Leakey	http://en.wikipedia.org/wiki/Louis_Leakey
Louis Lepke	http://en.wikipedia.org/wiki/Louis_Lepke
Louis MacNeice	http://en.wikipedia.org/wiki/Louis_MacNeice
Louis Malle	http://en.wikipedia.org/wiki/Louis_Malle
Louis McHenry Howe	http://en.wikipedia.org/wiki/Louis_McHenry_Howe
Louis Menand	http://en.wikipedia.org/wiki/Louis_Menand
Louis N�el	http://en.wikipedia.org/wiki/Louis_N%C3%A9el
Louis Nizer	http://en.wikipedia.org/wiki/Louis_Nizer
Louis Pasteur	http://en.wikipedia.org/wiki/Louis_Pasteur
Louis Philippe Joseph, duc d'Orl�ans	http://en.wikipedia.org/wiki/Louis_Philippe_Joseph,_duc_d%27Orl%C3%A9ans
Louis Renault	http://en.wikipedia.org/wiki/Louis_Renault_%28jurist%29
Louis Rukeyser	http://en.wikipedia.org/wiki/Louis_Rukeyser
Louis Simpson	http://en.wikipedia.org/wiki/Louis_Simpson
Louis St. Laurent	http://en.wikipedia.org/wiki/Louis_St._Laurent
Louis Stokes	http://en.wikipedia.org/wiki/Louis_Stokes
Louis Sullivan	http://en.wikipedia.org/wiki/Louis_Sullivan
Louis the Stammerer	http://en.wikipedia.org/wiki/Louis_the_Stammerer
Louis Theroux	http://en.wikipedia.org/wiki/Louis_Theroux
Louis Untermeyer	http://en.wikipedia.org/wiki/Louis_Untermeyer
Louis V	http://en.wikipedia.org/wiki/Louis_V_of_France
Louis V. Gerstner	http://en.wikipedia.org/wiki/Louis_V._Gerstner,_Jr.
Louis VI	http://en.wikipedia.org/wiki/Louis_VI_of_France
Louis VII	http://en.wikipedia.org/wiki/Louis_VII_of_France
Louis VIII	http://en.wikipedia.org/wiki/Louis_VIII_of_France
Louis Vuitton	http://en.wikipedia.org/wiki/Louis_Vuitton
Louis X	http://en.wikipedia.org/wiki/Louis_X_of_France
Louis XI	http://en.wikipedia.org/wiki/Louis_XI_of_France
Louis XII	http://en.wikipedia.org/wiki/Louis_XII_of_France
Louis XIII	http://en.wikipedia.org/wiki/Louis_XIII_of_France
Louis XIV	http://en.wikipedia.org/wiki/Louis_XIV_of_France
Louis XV	http://en.wikipedia.org/wiki/Louis_XV_of_France
Louis XVI	http://en.wikipedia.org/wiki/Louis_XVI_of_France
Louis XVII	http://en.wikipedia.org/wiki/Louis_XVII_of_France
Louis XVIII	http://en.wikipedia.org/wiki/Louis_XVIII_of_France
Louis Zukofsky	http://en.wikipedia.org/wiki/Louis_Zukofsky
Louisa May Alcott	http://en.wikipedia.org/wiki/Louisa_May_Alcott
Louise Bagshawe	http://en.wikipedia.org/wiki/Louise_Bagshawe
Louise Beavers	http://en.wikipedia.org/wiki/Louise_Beavers
Louise Bogan	http://en.wikipedia.org/wiki/Louise_Bogan
Louise Brooks	http://en.wikipedia.org/wiki/Louise_Brooks
Louise Ellman	http://en.wikipedia.org/wiki/Louise_Ellman
Louise Erdrich	http://en.wikipedia.org/wiki/Louise_Erdrich
Louise Fletcher	http://en.wikipedia.org/wiki/Louise_Fletcher
Louise Gl�ck	http://en.wikipedia.org/wiki/Louise_Gl%C3%BCck
Louise Imogen Guiney	http://en.wikipedia.org/wiki/Louise_Imogen_Guiney
Louise Jameson	http://en.wikipedia.org/wiki/Louise_Jameson
Louise Lasser	http://en.wikipedia.org/wiki/Louise_Lasser
Louise Mandrell	http://en.wikipedia.org/wiki/Louise_Mandrell
Louise Nevelson	http://en.wikipedia.org/wiki/Louise_Nevelson
Louise of Savoy	http://en.wikipedia.org/wiki/Louise_of_Savoy
Louise Post	http://en.wikipedia.org/wiki/Louise_Post
Louise Rainer	http://en.wikipedia.org/wiki/Louise_Rainer
Louise Slaughter	http://en.wikipedia.org/wiki/Louise_Slaughter
Louis-Ferdinand C�line	http://en.wikipedia.org/wiki/Louis-Ferdinand_C%C3%A9line
Louis-Jacques Th�nard	http://en.wikipedia.org/wiki/Louis_Jacques_Th%C3%A9nard
Louis-Jean-Marie Daubenton	http://en.wikipedia.org/wiki/Louis-Jean-Marie_Daubenton
Louis-Joseph, duc de Vend�me	http://en.wikipedia.org/wiki/Louis_Joseph,_duc_de_Vend%C3%B4me
Louis-Nicolas Davout	http://en.wikipedia.org/wiki/Louis-Nicolas_Davout
Lowell Bergman	http://en.wikipedia.org/wiki/Lowell_Bergman
Lowell Fulson	http://en.wikipedia.org/wiki/Lowell_Fulson
Lowell Jacoby	http://en.wikipedia.org/wiki/Lowell_E._Jacoby
Lowell P. Weicker, Jr.	http://en.wikipedia.org/wiki/Lowell_P._Weicker,_Jr.
Lowell Thomas	http://en.wikipedia.org/wiki/Lowell_Thomas
Luc Besson	http://en.wikipedia.org/wiki/Luc_Besson
Luc Holste	http://en.wikipedia.org/wiki/Luc_Holste
Luca Giordano	http://en.wikipedia.org/wiki/Luca_Giordano
Lucas Black	http://en.wikipedia.org/wiki/Lucas_Black
Lucas Cranach	http://en.wikipedia.org/wiki/Lucas_Cranach_the_Elder
Lucas van Leyden	http://en.wikipedia.org/wiki/Lucas_van_Leyden
Luchino Visconti	http://en.wikipedia.org/wiki/Luchino_Visconti
Luciana Berger	http://en.wikipedia.org/wiki/Luciana_Berger
Luciano Berio	http://en.wikipedia.org/wiki/Luciano_Berio
Luciano Pavarotti	http://en.wikipedia.org/wiki/Luciano_Pavarotti
Lucie Arnaz	http://en.wikipedia.org/wiki/Lucie_Arnaz
Lucien Ballard	http://en.wikipedia.org/wiki/Lucien_Ballard
Lucille Ball	http://en.wikipedia.org/wiki/Lucille_Ball
Lucille Bremer	http://en.wikipedia.org/wiki/Lucille_Bremer
Lucille Clifton	http://en.wikipedia.org/wiki/Lucille_Clifton
Lucille Roybal-Allard	http://en.wikipedia.org/wiki/Lucille_Roybal-Allard
Lucinda Williams	http://en.wikipedia.org/wiki/Lucinda_Williams
Lucine Amara	http://en.wikipedia.org/wiki/Lucine_Amara
Lucio Agostini	http://en.wikipedia.org/wiki/Lucio_Agostini
Lucius Licinius Lucullus	http://en.wikipedia.org/wiki/Lucius_Licinius_Lucullus
Lucius Verus	http://en.wikipedia.org/wiki/Lucius_Verus
Lucky Luciano	http://en.wikipedia.org/wiki/Lucky_Luciano
Lucretia Mott	http://en.wikipedia.org/wiki/Lucretia_Mott
Lucretia Peabody Hale	http://en.wikipedia.org/wiki/Lucretia_Peabody_Hale
Lucrezia Borgia	http://en.wikipedia.org/wiki/Lucrezia_Borgia
Lucy Briers	http://en.wikipedia.org/wiki/Lucy_Briers
Lucy Lawless	http://en.wikipedia.org/wiki/Lucy_Lawless
Lucy Liu	http://en.wikipedia.org/wiki/Lucy_Liu
Lucy Maud Montgomery	http://en.wikipedia.org/wiki/Lucy_Maud_Montgomery
Lucy Walter	http://en.wikipedia.org/wiki/Lucy_Walter
Ludivine Sagnier	http://en.wikipedia.org/wiki/Ludivine_Sagnier
Ludovic Hal�vy	http://en.wikipedia.org/wiki/Ludovic_Hal%e9vy
Ludovico Ariosto	http://en.wikipedia.org/wiki/Ludovico_Ariosto
Ludvig Holberg	http://en.wikipedia.org/wiki/Ludvig_Holberg
Ludwig Beck	http://en.wikipedia.org/wiki/Ludwig_Beck
Ludwig Berger	http://en.wikipedia.org/wiki/Ludwig_Berger_%28director%29
Ludwig Erhard	http://en.wikipedia.org/wiki/Ludwig_Erhard
Ludwig Feuerbach	http://en.wikipedia.org/wiki/Ludwig_Feuerbach
Ludwig Haetzer	http://en.wikipedia.org/wiki/Ludwig_Haetzer
Ludwig II	http://en.wikipedia.org/wiki/Ludwig_II
Ludwig Mies van der Rohe	http://en.wikipedia.org/wiki/Ludwig_Mies_van_der_Rohe
Ludwig Prandtl	http://en.wikipedia.org/wiki/Ludwig_Prandtl
Ludwig Quidde	http://en.wikipedia.org/wiki/Ludwig_Quidde
Ludwig Scotty	http://en.wikipedia.org/wiki/Ludwig_Scotty
Ludwig Tieck	http://en.wikipedia.org/wiki/Ludwig_Tieck
Ludwig van Beethoven	http://en.wikipedia.org/wiki/Ludwig_van_Beethoven
Ludwig von Mises	http://en.wikipedia.org/wiki/Ludwig_von_Mises
Ludwig Wittgenstein	http://en.wikipedia.org/wiki/Ludwig_Wittgenstein
Luigi Boccherini	http://en.wikipedia.org/wiki/Luigi_Boccherini
Luigi Cherubini	http://en.wikipedia.org/wiki/Luigi_Cherubini
Luigi Cornaro	http://en.wikipedia.org/wiki/Luigi_Cornaro
Luigi Dallapiccola	http://en.wikipedia.org/wiki/Luigi_Dallapiccola
Luigi Galvani	http://en.wikipedia.org/wiki/Luigi_Galvani
Luigi Nono	http://en.wikipedia.org/wiki/Luigi_Nono
Luigi Pirandello	http://en.wikipedia.org/wiki/Luigi_Pirandello
Luigi Russolo	http://en.wikipedia.org/wiki/Luigi_Russolo
Luis Alberni	http://en.wikipedia.org/wiki/Luis_Alberni
Luis Alfredo Garavito	http://en.wikipedia.org/wiki/Luis_Alfredo_Garavito
Luis Bu�uel	http://en.wikipedia.org/wiki/Luis_Bu%f1uel
Luis Cernuda	http://en.wikipedia.org/wiki/Luis_Cernuda
Lu�s de Cam�es	http://en.wikipedia.org/wiki/Lu%eds_de_Cam%f5es
Lu�s de G�ngora y Argote	http://en.wikipedia.org/wiki/Lu%eds_de_G%f3ngora_y_Argote
Luis Figo	http://en.wikipedia.org/wiki/Luis_Figo
Lu�s Figo	http://en.wikipedia.org/wiki/Lu%eds_Figo
Luis Fortuno	http://en.wikipedia.org/wiki/Luis_Fortuno
Luis Gutierrez	http://en.wikipedia.org/wiki/Luis_Gutierrez
Luis Guzm�n	http://en.wikipedia.org/wiki/Luis_Guzm%e1n
Luis Leloir	http://en.wikipedia.org/wiki/Luis_Leloir
Luis Miguel	http://en.wikipedia.org/wiki/Luis_Miguel
Luis Pal�s Matos	http://en.wikipedia.org/wiki/Luis_Pal%e9s_Matos
Luis Posada Carriles	http://en.wikipedia.org/wiki/Luis_Posada_Carriles
Luis W. Alvarez	http://en.wikipedia.org/wiki/Luis_W._Alvarez
Luisa Diogo	http://en.wikipedia.org/wiki/Luisa_Diogo
Luisa Diogo	http://en.wikipedia.org/wiki/Luisa_Diogo
Luiz In�cio Lula da Silva	http://en.wikipedia.org/wiki/Luiz_In%e1cio_Lula_da_Silva
Lukas Haas	http://en.wikipedia.org/wiki/Lukas_Haas
Luke Ford	http://en.wikipedia.org/wiki/Luke_Ford
Luke Halpin	http://en.wikipedia.org/wiki/Luke_Halpin
Luke Hansard	http://en.wikipedia.org/wiki/Luke_Hansard
Luke Perry	http://en.wikipedia.org/wiki/Luke_Perry
Luke Vibert	http://en.wikipedia.org/wiki/Luke_Vibert
Luke Wilson	http://en.wikipedia.org/wiki/Luke_Wilson
Lung Leg	http://en.wikipedia.org/wiki/Lung_Leg
Lupe Velez	http://en.wikipedia.org/wiki/Lupe_Velez
Lurleen Burns Wallace	http://en.wikipedia.org/wiki/Lurleen_Burns_Wallace
Luther Allison	http://en.wikipedia.org/wiki/Luther_Allison
Luther Burbank	http://en.wikipedia.org/wiki/Luther_Burbank
Luther Campbell	http://en.wikipedia.org/wiki/Luther_Campbell
Luther Vandross	http://en.wikipedia.org/wiki/Luther_Vandross
Lutz Schwerin von Krosigk	http://en.wikipedia.org/wiki/Lutz_Schwerin_von_Krosigk
Lydia Lunch	http://en.wikipedia.org/wiki/Lydia_Lunch
Lyle Alzado	http://en.wikipedia.org/wiki/Lyle_Alzado
Lyle Alzado	http://en.wikipedia.org/wiki/Lyle_Alzado
Lyle Lovett	http://en.wikipedia.org/wiki/Lyle_Lovett
Lyle Menendez	http://en.wikipedia.org/wiki/Lyle_Menendez
Lyle Talbot	http://en.wikipedia.org/wiki/Lyle_Talbot
Lyle Waggoner	http://en.wikipedia.org/wiki/Lyle_Waggoner
Lyman Beecher	http://en.wikipedia.org/wiki/Lyman_Beecher
Lyman Knapp	http://en.wikipedia.org/wiki/Lyman_Knapp
Lyn Brown	http://en.wikipedia.org/wiki/Lyn_Brown_%28journalist%29
Lyn Collins	http://en.wikipedia.org/wiki/Lyn_Collins
Lyn Nofziger	http://en.wikipedia.org/wiki/Lyn_Nofziger
Lynd Ward	http://en.wikipedia.org/wiki/Lynd_Ward
Lynda Barry	http://en.wikipedia.org/wiki/Lynda_Barry
Lynda Carter	http://en.wikipedia.org/wiki/Lynda_Carter
Lynda Day George	http://en.wikipedia.org/wiki/Lynda_Day_George
Lynden Oscar Pindling	http://en.wikipedia.org/wiki/Lynden_Oscar_Pindling
Lyndon B. Johnson	http://en.wikipedia.org/wiki/Lyndon_B._Johnson
Lyndon LaRouche	http://en.wikipedia.org/wiki/Lyndon_LaRouche
Lynn Abbey	http://en.wikipedia.org/wiki/Lynn_Abbey
Lynn Anderson	http://en.wikipedia.org/wiki/Lynn_Anderson
Lynn Bari	http://en.wikipedia.org/wiki/Lynn_Bari
Lynn Fontanne	http://en.wikipedia.org/wiki/Lynn_Fontanne
Lynn Jenkins	http://en.wikipedia.org/wiki/Lynn_Jenkins
Lynn Johnston	http://en.wikipedia.org/wiki/Lynn_Johnston
Lynn Martin	http://en.wikipedia.org/wiki/Lynn_Martin
Lynn Martin	http://en.wikipedia.org/wiki/Lynn_Martin
Lynn Redgrave	http://en.wikipedia.org/wiki/Lynn_Redgrave
Lynn Swann	http://en.wikipedia.org/wiki/Lynn_Swann
Lynn Westmoreland	http://en.wikipedia.org/wiki/Lynn_Westmoreland
Lynn Whitfield	http://en.wikipedia.org/wiki/Lynn_Whitfield
Lynn Woolsey	http://en.wikipedia.org/wiki/Lynn_Woolsey
Lynndie England	http://en.wikipedia.org/wiki/Lynndie_England
Lynne Cheney	http://en.wikipedia.org/wiki/Lynne_Cheney
Lynne Featherstone	http://en.wikipedia.org/wiki/Lynne_Featherstone
Lynne Ramsay	http://en.wikipedia.org/wiki/Lynne_Ramsay
Lynne Thigpen	http://en.wikipedia.org/wiki/Lynne_Thigpen
Lynx Gaede	http://en.wikipedia.org/wiki/Lynx_Gaede
Lyonpo Sangay Ngedup	http://en.wikipedia.org/wiki/Lyonpo_Sangay_Ngedup
Lytton Strachey	http://en.wikipedia.org/wiki/Lytton_Strachey
M. C. Escher	http://en.wikipedia.org/wiki/M._C._Escher
M. Emmet Walsh	http://en.wikipedia.org/wiki/M._Emmet_Walsh
M. Jodi Rell	http://en.wikipedia.org/wiki/M._Jodi_Rell
M. Night Shyamalan	http://en.wikipedia.org/wiki/M._Night_Shyamalan
M. R. James	http://en.wikipedia.org/wiki/M._R._James
M. Scott Peck	http://en.wikipedia.org/wiki/M._Scott_Peck
Ma Barker	http://en.wikipedia.org/wiki/Ma_Barker
Ma Ying-jeou	http://en.wikipedia.org/wiki/Ma_Ying-jeou
Maatia Toafa	http://en.wikipedia.org/wiki/Maatia_Toafa
Mabel Dodge Luhan	http://en.wikipedia.org/wiki/Mabel_Dodge_Luhan
Mabel King	http://en.wikipedia.org/wiki/Mabel_King
Mabel Normand	http://en.wikipedia.org/wiki/Mabel_Normand
Mac Bundy	http://en.wikipedia.org/wiki/Mac_Bundy
Mac Collins	http://en.wikipedia.org/wiki/Mac_Collins
Mac Davis	http://en.wikipedia.org/wiki/Mac_Davis
Mac Dre	http://en.wikipedia.org/wiki/Mac_Dre
Mac Sweeney	http://en.wikipedia.org/wiki/Mac_Sweeney
Mac Thornberry	http://en.wikipedia.org/wiki/Mac_Thornberry
Macaulay Culkin	http://en.wikipedia.org/wiki/Macaulay_Culkin
Macedonio Melloni	http://en.wikipedia.org/wiki/Macedonio_Melloni
Machado de Assis	http://en.wikipedia.org/wiki/Machado_de_Assis
Mack 10	http://en.wikipedia.org/wiki/Mack_10
Mack Mattingly	http://en.wikipedia.org/wiki/Mack_Mattingly
Mack McLarty	http://en.wikipedia.org/wiki/Mack_McLarty
Mack Sennett	http://en.wikipedia.org/wiki/Mack_Sennett
Mackenzie Astin	http://en.wikipedia.org/wiki/Mackenzie_Astin
Mackenzie Bowell	http://en.wikipedia.org/wiki/Mackenzie_Bowell
Mackenzie Crook	http://en.wikipedia.org/wiki/Mackenzie_Crook
Mackenzie Phillips	http://en.wikipedia.org/wiki/Mackenzie_Phillips
Mackenzie Rosman	http://en.wikipedia.org/wiki/Mackenzie_Rosman
MacKinlay Kantor	http://en.wikipedia.org/wiki/MacKinlay_Kantor
Macky Sall	http://en.wikipedia.org/wiki/Macky_Sall
Macy Gray	http://en.wikipedia.org/wiki/Macy_Gray
Madalyn Murray O'Hair	http://en.wikipedia.org/wiki/Madalyn_Murray_O'Hair
Madame Chiang Kai-Shek	http://en.wikipedia.org/wiki/Madame_Chiang_Kai-Shek
Madame de S�vign�	http://en.wikipedia.org/wiki/Madame_de_S%e9vign%e9
Madame de Sta�l	http://en.wikipedia.org/wiki/Madame_de_Sta%ebl
Madame Tussaud	http://en.wikipedia.org/wiki/Madame_Tussaud
M�dchen Amick	http://en.wikipedia.org/wiki/M%E4dchen_Amick
Madeleine Albright	http://en.wikipedia.org/wiki/Madeleine_Albright
Madeleine Bordallo	http://en.wikipedia.org/wiki/Madeleine_Bordallo
Madeleine Carroll	http://en.wikipedia.org/wiki/Madeleine_Carroll
Madeleine L'Engle	http://en.wikipedia.org/wiki/Madeleine_L'Engle
Madeleine Moon	http://en.wikipedia.org/wiki/Madeleine_Moon
Madeleine Stowe	http://en.wikipedia.org/wiki/Madeleine_Stowe
Madeline Kahn	http://en.wikipedia.org/wiki/Madeline_Kahn
Madeline Zima	http://en.wikipedia.org/wiki/Madeline_Zima
Madge Evans	http://en.wikipedia.org/wiki/Madge_Evans
Madhav Kumar Nepal	http://en.wikipedia.org/wiki/Madhav_Kumar_Nepal
Mae Murray	http://en.wikipedia.org/wiki/Mae_Murray
Mae West	http://en.wikipedia.org/wiki/Mae_West
Mae Whitman	http://en.wikipedia.org/wiki/Mae_Whitman
M�rsk Mc-Kinney M�ller	http://en.wikipedia.org/wiki/M%E6rsk_Mc-Kinney_M%F8ller
Magali Amadei	http://en.wikipedia.org/wiki/Magali_Amadei
Magda Gabor	http://en.wikipedia.org/wiki/Magda_Gabor
Magdalena Wrobel	http://en.wikipedia.org/wiki/Magdalena_Wrobel
Maggie Grace	http://en.wikipedia.org/wiki/Maggie_Grace
Maggie Gyllenhaal	http://en.wikipedia.org/wiki/Maggie_Gyllenhaal
Maggie Kuhn	http://en.wikipedia.org/wiki/Maggie_Kuhn
Maggie Smith	http://en.wikipedia.org/wiki/Maggie_Smith
Magic Johnson	http://en.wikipedia.org/wiki/Magic_Johnson
Mahalia Jackson	http://en.wikipedia.org/wiki/Mahalia_Jackson
Mahamadou Danda	http://en.wikipedia.org/wiki/Mahamadou_Danda
Maharishi Mahesh Yogi	http://en.wikipedia.org/wiki/Maharishi_Mahesh_Yogi
Mahatma Gandhi	http://en.wikipedia.org/wiki/Mahatma_Gandhi
Mahendra Singh Dhoni	http://en.wikipedia.org/wiki/Mahendra_Singh_Dhoni
Mahinda Rajapakse	http://en.wikipedia.org/wiki/Mahinda_Rajapakse
Mahmood Mamdani	http://en.wikipedia.org/wiki/Mahmood_Mamdani
Mahmoud Abbas	http://en.wikipedia.org/wiki/Mahmoud_Abbas
Mahmoud Ahmad	http://en.wikipedia.org/wiki/Mahmoud_Ahmad
Mahmoud Ahmadinejad	http://en.wikipedia.org/wiki/Mahmoud_Ahmadinejad
Mahmoud Zahar	http://en.wikipedia.org/wiki/Mahmoud_Zahar
Mairead Corrigan	http://en.wikipedia.org/wiki/Mairead_Corrigan
Majel Barrett	http://en.wikipedia.org/wiki/Majel_Barrett
Major Owens	http://en.wikipedia.org/wiki/Major_Owens
Maktoum bin Rashid al-Maktoum	http://en.wikipedia.org/wiki/Maktoum_bin_Rashid_al-Maktoum
Malachi Favors	http://en.wikipedia.org/wiki/Malachi_Favors
Malachi York-El	http://en.wikipedia.org/wiki/Malachi_York-El
Malachy McCourt	http://en.wikipedia.org/wiki/Malachy_McCourt
Malam Bacai Sanh�	http://en.wikipedia.org/wiki/Malam_Bacai_Sanh%E1
Malcolm Baldrige	http://en.wikipedia.org/wiki/Malcolm_Baldrige,_Jr.
Malcolm Bradbury	http://en.wikipedia.org/wiki/Malcolm_Bradbury
Malcolm Bruce	http://en.wikipedia.org/wiki/Malcolm_Bruce
Malcolm Cowley	http://en.wikipedia.org/wiki/Malcolm_Cowley
Malcolm David Kelley	http://en.wikipedia.org/wiki/Malcolm_David_Kelley
Malcolm Forbes	http://en.wikipedia.org/wiki/Malcolm_Forbes
Malcolm Fraser	http://en.wikipedia.org/wiki/Malcolm_Fraser
Malcolm Gladwell	http://en.wikipedia.org/wiki/Malcolm_Gladwell
Malcolm Lowry	http://en.wikipedia.org/wiki/Malcolm_Lowry
Malcolm Marshall	http://en.wikipedia.org/wiki/Malcolm_Marshall
Malcolm McDowell	http://en.wikipedia.org/wiki/Malcolm_McDowell
Malcolm McLaren	http://en.wikipedia.org/wiki/Malcolm_McLaren
Malcolm Muggeridge	http://en.wikipedia.org/wiki/Malcolm_Muggeridge
Malcolm Rifkind	http://en.wikipedia.org/wiki/Malcolm_Rifkind
Malcolm Wallop	http://en.wikipedia.org/wiki/Malcolm_Wallop
Malcolm Wicks	http://en.wikipedia.org/wiki/Malcolm_Wicks
Malcolm Wilson	http://en.wikipedia.org/wiki/Malcolm_Wilson_(governor)
Malcolm X	http://en.wikipedia.org/wiki/Malcolm_X
Malcolm Young	http://en.wikipedia.org/wiki/Malcolm_Young
Malcolm-Jamal Warner	http://en.wikipedia.org/wiki/Malcolm-Jamal_Warner
Malietoa Tanumafili II	http://en.wikipedia.org/wiki/Malietoa_Tanumafili_II
Malin Akerman	http://en.wikipedia.org/wiki/Malin_Akerman
Malinda Williams	http://en.wikipedia.org/wiki/Malinda_Williams
Mama Cass	http://en.wikipedia.org/wiki/Mama_Cass
Mamie Eisenhower	http://en.wikipedia.org/wiki/Mamie_Eisenhower
Mamie Van Doren	http://en.wikipedia.org/wiki/Mamie_Van_Doren
Man Ray	http://en.wikipedia.org/wiki/Man_Ray
Manasseh Sogavare	http://en.wikipedia.org/wiki/Manasseh_Sogavare
Mandy Moore	http://en.wikipedia.org/wiki/Mandy_Moore
Mandy Patinkin	http://en.wikipedia.org/wiki/Mandy_Patinkin
Manfred Eigen	http://en.wikipedia.org/wiki/Manfred_Eigen
Manfred Mann	http://en.wikipedia.org/wiki/Manfred_Mann_(musician)
Mangosuthu Buthelezi	http://en.wikipedia.org/wiki/Mangosuthu_Buthelezi
Manmohan Singh	http://en.wikipedia.org/wiki/Manmohan_Singh
Manne Siegbahn	http://en.wikipedia.org/wiki/Manne_Siegbahn
Mannie Fresh	http://en.wikipedia.org/wiki/Mannie_Fresh
Manny Alvarez	http://en.wikipedia.org/wiki/Manny_Alvarez
Manny Mori	http://en.wikipedia.org/wiki/Manny_Mori
Manny Ramirez	http://en.wikipedia.org/wiki/Manny_Ramirez
Manuel de Falla	http://en.wikipedia.org/wiki/Manuel_de_Falla
Manuel I Comnenus	http://en.wikipedia.org/wiki/Manuel_I_Comnenus
Manuel II Palaeologus	http://en.wikipedia.org/wiki/Manuel_II_Palaeologus
Manuel Lujan, Jr.	http://en.wikipedia.org/wiki/Manuel_Lujan%2C_Jr.
Manuel Noriega	http://en.wikipedia.org/wiki/Manuel_Noriega
Manuel Philes	http://en.wikipedia.org/wiki/Manuel_Philes
Manuel Puig	http://en.wikipedia.org/wiki/Manuel_Puig
Manuel Quezon	http://en.wikipedia.org/wiki/Manuel_Quezon
Manuel Roxas	http://en.wikipedia.org/wiki/Manuel_Roxas
Manuel Tamayo y Baus	http://en.wikipedia.org/wiki/Manuel_Tamayo_y_Baus
Manuel Zelaya	http://en.wikipedia.org/wiki/Manuel_Zelaya
Manute Bol	http://en.wikipedia.org/wiki/Manute_Bol
Mara Corday	http://en.wikipedia.org/wiki/Mara_Corday
Mara Liasson	http://en.wikipedia.org/wiki/Mara_Liasson
Mara Wilson	http://en.wikipedia.org/wiki/Mara_Wilson
Marat Safin	http://en.wikipedia.org/wiki/Marat_Safin
Marc Alfos	http://en.wikipedia.org/wiki/Marc_Alfos
Marc All�gret	http://en.wikipedia.org/wiki/Marc_All%E9gret
Marc Almond	http://en.wikipedia.org/wiki/Marc_Almond
Marc Andreessen	http://en.wikipedia.org/wiki/Marc_Andreessen
Marc Anthony	http://en.wikipedia.org/wiki/Marc_Anthony
Marc Blank	http://en.wikipedia.org/wiki/Marc_Blank
Marc Blitzstein	http://en.wikipedia.org/wiki/Marc_Blitzstein
Marc Blucas	http://en.wikipedia.org/wiki/Marc_Blucas
Marc Bolan	http://en.wikipedia.org/wiki/Marc_Bolan
Marc Chagall	http://en.wikipedia.org/wiki/Marc_Chagall
Marc Cohn	http://en.wikipedia.org/wiki/Marc_Cohn
Marc Dutroux	http://en.wikipedia.org/wiki/Marc_Dutroux
Marc Jacobs	http://en.wikipedia.org/wiki/Marc_Jacobs
Marc Klaas	http://en.wikipedia.org/wiki/Marc_Klaas
Marc Lawrence	http://en.wikipedia.org/wiki/Marc_Lawrence
Marc Maron	http://en.wikipedia.org/wiki/Marc_Maron
Marc Morial	http://en.wikipedia.org/wiki/Marc_Morial
Marc Racicot	http://en.wikipedia.org/wiki/Marc_Racicot
Marc Ravalomanana	http://en.wikipedia.org/wiki/Marc_Ravalomanana
Marc Ribot	http://en.wikipedia.org/wiki/Marc_Ribot
Marc Rich	http://en.wikipedia.org/wiki/Marc_Rich
Marc Rotenberg	http://en.wikipedia.org/wiki/Marc_Rotenberg
Marc Singer	http://en.wikipedia.org/wiki/Marc_Singer
Marcel Breuer	http://en.wikipedia.org/wiki/Marcel_Breuer
Marcel Carn�	http://en.wikipedia.org/wiki/Marcel_Carn%E9
Marcel Duchamp	http://en.wikipedia.org/wiki/Marcel_Duchamp
Marcel Dupr�	http://en.wikipedia.org/wiki/Marcel_Dupr%E9
Marcel Marceau	http://en.wikipedia.org/wiki/Marcel_Marceau
Marcel Mauss	http://en.wikipedia.org/wiki/Marcel_Mauss
Marcel Proust	http://en.wikipedia.org/wiki/Marcel_Proust
Marcellin Berthelot	http://en.wikipedia.org/wiki/Marcellin_Berthelot
Marcello Abbado	http://en.wikipedia.org/wiki/Marcello_Abbado
Marcello Malpighi	http://en.wikipedia.org/wiki/Marcello_Malpighi
Marcello Mastroianni	http://en.wikipedia.org/wiki/Marcello_Mastroianni
Marcello Mastroianni	http://en.wikipedia.org/wiki/Marcello_Mastroianni
Marcia C. Kaptur	http://en.wikipedia.org/wiki/Marcia_C._Kaptur
Marcia Cross	http://en.wikipedia.org/wiki/Marcia_Cross
Marcia Fudge	http://en.wikipedia.org/wiki/Marcia_Fudge
Marcia Gay Harden	http://en.wikipedia.org/wiki/Marcia_Gay_Harden
Marcia Wallace	http://en.wikipedia.org/wiki/Marcia_Wallace
Marco Conti	http://en.wikipedia.org/wiki/Marco_Conti
Marco Polo	http://en.wikipedia.org/wiki/Marco_Polo
Marco van Basten	http://en.wikipedia.org/wiki/Marco_van_Basten
Marcus Allen	http://en.wikipedia.org/wiki/Marcus_Allen
Marcus Alonzo Hanna	http://en.wikipedia.org/wiki/Marcus_Alonzo_Hanna
Marcus Aurelius	http://en.wikipedia.org/wiki/Marcus_Aurelius
Marcus Camby	http://en.wikipedia.org/wiki/Marcus_Camby
Marcus Garvey	http://en.wikipedia.org/wiki/Marcus_Garvey
Marcus Jones	http://en.wikipedia.org/wiki/Marcus_Jones_(UK_politician)
Marcus Schenkenberg	http://en.wikipedia.org/wiki/Marcus_Schenkenberg
Marcus Stephen	http://en.wikipedia.org/wiki/Marcus_Stephen
Marcy Kaptur	http://en.wikipedia.org/wiki/Marcy_Kaptur
Mare Winningham	http://en.wikipedia.org/wiki/Mare_Winningham
Marek Belka	http://en.wikipedia.org/wiki/Marek_Belka
Marg Helgenberger	http://en.wikipedia.org/wiki/Marg_Helgenberger
Margaret Anderson	http://en.wikipedia.org/wiki/Margaret_Anderson
Margaret Atwood	http://en.wikipedia.org/wiki/Margaret_Atwood
Margaret Beckett	http://en.wikipedia.org/wiki/Margaret_Beckett
Margaret Booth	http://en.wikipedia.org/wiki/Margaret_Booth
Margaret Carlson	http://en.wikipedia.org/wiki/Margaret_Carlson
Margaret Chase Smith	http://en.wikipedia.org/wiki/Margaret_Chase_Smith
Margaret Cho	http://en.wikipedia.org/wiki/Margaret_Cho
Margaret Curran	http://en.wikipedia.org/wiki/Margaret_Curran
Margaret Deland	http://en.wikipedia.org/wiki/Margaret_Deland
Margaret Drabble	http://en.wikipedia.org/wiki/Margaret_Drabble
Margaret Dumont	http://en.wikipedia.org/wiki/Margaret_Dumont
Margaret Fuller	http://en.wikipedia.org/wiki/Margaret_Fuller
Margaret Hamilton	http://en.wikipedia.org/wiki/Margaret_Hamilton
Margaret Hayes	http://en.wikipedia.org/wiki/Margaret_Hayes
Margaret Hodge	http://en.wikipedia.org/wiki/Margaret_Hodge
Margaret Kennedy	http://en.wikipedia.org/wiki/Margaret_Kennedy
Margaret Leighton	http://en.wikipedia.org/wiki/Margaret_Leighton
Margaret Lockwood	http://en.wikipedia.org/wiki/Margaret_Lockwood
Margaret Mead	http://en.wikipedia.org/wiki/Margaret_Mead
Margaret Mitchell	http://en.wikipedia.org/wiki/Margaret_Mitchell
Margaret Murray	http://en.wikipedia.org/wiki/Margaret_Murray
Margaret O'Brien	http://en.wikipedia.org/wiki/Margaret_O%27Brien
Margaret of Angoul�me	http://en.wikipedia.org/wiki/Margaret_of_Angoul%EAme
Margaret of Anjou	http://en.wikipedia.org/wiki/Margaret_of_Anjou
Margaret of Austria	http://en.wikipedia.org/wiki/Archduchess_Margarethe_Klementine_of_Austria
Margaret of Parma	http://en.wikipedia.org/wiki/Margaret_of_Parma
Margaret of Valois	http://en.wikipedia.org/wiki/Margaret_of_Valois
Margaret Oliphant	http://en.wikipedia.org/wiki/Margaret_Oliphant
Margaret O'Neill Eaton	http://en.wikipedia.org/wiki/Margaret_O%27Neill_Eaton
Margaret Peterson Haddix	http://en.wikipedia.org/wiki/Margaret_Peterson_Haddix
Margaret Ritchie	http://en.wikipedia.org/wiki/Margaret_Ritchie_(politician)
Margaret Rutherford	http://en.wikipedia.org/wiki/Margaret_Rutherford
Margaret Sanger	http://en.wikipedia.org/wiki/Margaret_Sanger
Margaret Spellings	http://en.wikipedia.org/wiki/Margaret_Spellings
Margaret Thatcher	http://en.wikipedia.org/wiki/Margaret_Thatcher
Margaret Truman	http://en.wikipedia.org/wiki/Margaret_Truman
Margaret Tudor	http://en.wikipedia.org/wiki/Margaret_Tudor
Margaret Walker	http://en.wikipedia.org/wiki/Margaret_Walker
Margaux Hemingway	http://en.wikipedia.org/wiki/Margaux_Hemingway
Marge Piercy	http://en.wikipedia.org/wiki/Marge_Piercy
Marge Roukema	http://en.wikipedia.org/wiki/Marge_Roukema
Marge Roukema	http://en.wikipedia.org/wiki/Marge_Roukema
Marge Schott	http://en.wikipedia.org/wiki/Marge_Schott
Margery Allingham	http://en.wikipedia.org/wiki/Margery_Allingham
Margi Clarke	http://en.wikipedia.org/wiki/Margi_Clarke
Margot Fonteyn	http://en.wikipedia.org/wiki/Margot_Fonteyn
Margot James	http://en.wikipedia.org/wiki/Margot_James
Margot Kidder	http://en.wikipedia.org/wiki/Margot_Kidder
Margrethe I	http://en.wikipedia.org/wiki/Margrethe_I
Margrethe II	http://en.wikipedia.org/wiki/Margrethe_II
Margrethe II	http://en.wikipedia.org/wiki/Margrethe_II
Marguerite Chapman	http://en.wikipedia.org/wiki/Marguerite_Chapman
Marguerite Duras	http://en.wikipedia.org/wiki/Marguerite_Duras
Marguerite Moreau	http://en.wikipedia.org/wiki/Marguerite_Moreau
Marguerite Young	http://en.wikipedia.org/wiki/Marguerite_Young
Marguerite Yourcenar	http://en.wikipedia.org/wiki/Marguerite_Yourcenar
Mar� Alkatiri	http://en.wikipedia.org/wiki/Mar%ED_Alkatiri
Mari Sandoz	http://en.wikipedia.org/wiki/Mari_Sandoz
Maria Bartiromo	http://en.wikipedia.org/wiki/Maria_Bartiromo
Maria Bello	http://en.wikipedia.org/wiki/Maria_Bello
Maria Callas	http://en.wikipedia.org/wiki/Maria_Callas
Maria Cantwell	http://en.wikipedia.org/wiki/Maria_Cantwell
Maria Conchita Alonso	http://en.wikipedia.org/wiki/Maria_Conchita_Alonso
Maria do Carmo Silveira	http://en.wikipedia.org/wiki/Maria_do_Carmo_Silveira
Maria Eagle	http://en.wikipedia.org/wiki/Maria_Eagle
Maria Edgeworth	http://en.wikipedia.org/wiki/Maria_Edgeworth
Maria Felix	http://en.wikipedia.org/wiki/Maria_Felix
Maria Gaetana Agnesi	http://en.wikipedia.org/wiki/Maria_Gaetana_Agnesi
Maria Goeppert-Mayer	http://en.wikipedia.org/wiki/Maria_Goeppert-Mayer
Maria Hinojosa	http://en.wikipedia.org/wiki/Maria_Hinojosa
Maria Innocentia Hummel	http://en.wikipedia.org/wiki/Maria_Innocentia_Hummel
Maria Menounos	http://en.wikipedia.org/wiki/Maria_Menounos
Maria Miller	http://en.wikipedia.org/wiki/Maria_Miller
Maria Montessori	http://en.wikipedia.org/wiki/Maria_Montessori
Maria Sharapova	http://en.wikipedia.org/wiki/Maria_Sharapova
Maria Shriver	http://en.wikipedia.org/wiki/Maria_Shriver
Maria Tallchief	http://en.wikipedia.org/wiki/Maria_Tallchief
Maria Theresa	http://en.wikipedia.org/wiki/Maria_Theresa
Mariah Carey	http://en.wikipedia.org/wiki/Mariah_Carey
Marian Anderson	http://en.wikipedia.org/wiki/Marian_Anderson
Marian Wright Edelman	http://en.wikipedia.org/wiki/Marian_Wright_Edelman
Mariann Aalda	http://en.wikipedia.org/wiki/Mariann_Aalda
Marianne Denicourt	http://en.wikipedia.org/wiki/Marianne_Denicourt
Marianne Faithfull	http://en.wikipedia.org/wiki/Marianne_Faithfull
Marianne Jean-Baptiste	http://en.wikipedia.org/wiki/Marianne_Jean-Baptiste
Marianne Moore	http://en.wikipedia.org/wiki/Marianne_Moore
Marie Am�lie Th�r�se	http://en.wikipedia.org/wiki/Maria_Amalia_of_Naples_and_Sicily
Marie Antoinette	http://en.wikipedia.org/wiki/Marie_Antoinette
Marie Blake	http://en.wikipedia.org/wiki/Marie_Blake
Marie Curie	http://en.wikipedia.org/wiki/Marie_Curie
Marie de France	http://en.wikipedia.org/wiki/Marie_de_France
Marie de Medici	http://en.wikipedia.org/wiki/Marie_de_Medici
Marie Dionne	http://en.wikipedia.org/wiki/Marie_Dionne
Marie Dressler	http://en.wikipedia.org/wiki/Marie_Dressler
Marie Leszczynska	http://en.wikipedia.org/wiki/Marie_Leszczynska
Marie Louise	http://en.wikipedia.org/wiki/Marie_Louise,_Duchess_of_Parma
Marie Osmond	http://en.wikipedia.org/wiki/Marie_Osmond
Marie Stopes	http://en.wikipedia.org/wiki/Marie_Stopes
Marie Th�r�se	http://en.wikipedia.org/wiki/Maria_Theresa_of_Spain
Marie Trintignant	http://en.wikipedia.org/wiki/Marie_Trintignant
Marie Wilson	http://en.wikipedia.org/wiki/Marie_Wilson_(American_actress)
Marie Windsor	http://en.wikipedia.org/wiki/Marie_Windsor
Marie-Fran�ois-Xavier Bichat	http://en.wikipedia.org/wiki/Marie_François_Xavier_Bichat
Mariel Hemingway	http://en.wikipedia.org/wiki/Mariel_Hemingway
Marie-No�lle Th�mereau	http://en.wikipedia.org/wiki/Marie-No%EBlle_Th%E9mereau
Mariette Hartley	http://en.wikipedia.org/wiki/Mariette_Hartley
Marilu Henner	http://en.wikipedia.org/wiki/Marilu_Henner
Marilyn Hacker	http://en.wikipedia.org/wiki/Marilyn_Hacker
Marilyn Horne	http://en.wikipedia.org/wiki/Marilyn_Horne
Marilyn Lloyd	http://en.wikipedia.org/wiki/Marilyn_Lloyd
Marilyn Manson	http://en.wikipedia.org/wiki/Marilyn_Manson
Marilyn Maxwell	http://en.wikipedia.org/wiki/Marilyn_Maxwell
Marilyn Monroe	http://en.wikipedia.org/wiki/Marilyn_Monroe
Marilyn Musgrave	http://en.wikipedia.org/wiki/Marilyn_Musgrave
Marilyn Quayle	http://en.wikipedia.org/wiki/Marilyn_Quayle
Marilyn vos Savant	http://en.wikipedia.org/wiki/Marilyn_vos_Savant
Marilyn Ware	http://en.wikipedia.org/wiki/Marilyn_Ware
Marilynne Robinson	http://en.wikipedia.org/wiki/Marilynne_Robinson
Marin Mersenne	http://en.wikipedia.org/wiki/Marin_Mersenne
Marina Sirtis	http://en.wikipedia.org/wiki/Marina_Sirtis
Marino Marini	http://en.wikipedia.org/wiki/Marino_Marini_(musician)
Mario Adorf	http://en.wikipedia.org/wiki/Mario_Adorf
Mario Andretti	http://en.wikipedia.org/wiki/Mario_Andretti
Mario Batali	http://en.wikipedia.org/wiki/Mario_Batali
Mario Biaggi	http://en.wikipedia.org/wiki/Mario_Biaggi
Mario Cantone	http://en.wikipedia.org/wiki/Mario_Cantone
Mario Cuomo	http://en.wikipedia.org/wiki/Mario_Cuomo
M�rio de S�-Carneiro	http://en.wikipedia.org/wiki/M%E1rio_de_S%E1-Carneiro
Mario Diaz-Balart	http://en.wikipedia.org/wiki/Mario_Diaz-Balart
Mario Gallo	http://en.wikipedia.org/wiki/Mario_Gallo_%28actor%29
Mario J. Molina	http://en.wikipedia.org/wiki/Mario_J._Molina
Mario Lanza	http://en.wikipedia.org/wiki/Mario_Lanza
Mario Lemieux	http://en.wikipedia.org/wiki/Mario_Lemieux
Mario Lopez	http://en.wikipedia.org/wiki/Mario_Lopez
Mario Monti	http://en.wikipedia.org/wiki/Mario_Monti
Mario Puzo	http://en.wikipedia.org/wiki/Mario_Puzo
M�rio Soares	http://en.wikipedia.org/wiki/M%E1rio_Soares
Mario Van Peebles	http://en.wikipedia.org/wiki/Mario_Van_Peebles
Mario Vargas Llosa	http://en.wikipedia.org/wiki/Mario_Vargas_Llosa
Marion Barry	http://en.wikipedia.org/wiki/Marion_Barry
Marion Berry	http://en.wikipedia.org/wiki/Robert_Marion_Berry
Marion Davies	http://en.wikipedia.org/wiki/Marion_Davies
Marion Jones	http://en.wikipedia.org/wiki/Marion_Jones
Marion Ross	http://en.wikipedia.org/wiki/Marion_Ross
Marion Zimmer Bradley	http://en.wikipedia.org/wiki/Marion_Zimmer_Bradley
Marisa Tomei	http://en.wikipedia.org/wiki/Marisa_Tomei
Mariska Hargitay	http://en.wikipedia.org/wiki/Mariska_Hargitay
Marjorie Courtenay-Latimer	http://en.wikipedia.org/wiki/Marjorie_Courtenay-Latimer
Marjorie Kinnan Rawlings	http://en.wikipedia.org/wiki/Marjorie_Kinnan_Rawlings
Marjorie Main	http://en.wikipedia.org/wiki/Marjorie_Main
Marjorie Rambeau	http://en.wikipedia.org/wiki/Marjorie_Rambeau
Marjorie S. Holt	http://en.wikipedia.org/wiki/Marjorie_S._Holt
Mark "Gator" Rogowski	http://en.wikipedia.org/wiki/Mark_Rogowski
Mark A. Altman	http://en.wikipedia.org/wiki/Mark_A._Altman
Mark Abene	http://en.wikipedia.org/wiki/Mark_Abene
Mark Addison	http://en.wikipedia.org/wiki/Mark_Addison
Mark Addy	http://en.wikipedia.org/wiki/Mark_Addy
Mark Amin	http://en.wikipedia.org/wiki/Mark_Amin
Mark Andrews	http://en.wikipedia.org/wiki/Mark_Andrews
Mark Antony	http://en.wikipedia.org/wiki/Mark_Antony
Mark Archer	http://en.wikipedia.org/wiki/Mark_Archer
Mark Begich	http://en.wikipedia.org/wiki/Mark_Begich
Mark Boucher	http://en.wikipedia.org/wiki/Mark_Boucher
Mark Burnett	http://en.wikipedia.org/wiki/Mark_Burnett
Mark C. Pigott	http://en.wikipedia.org/wiki/Mark_Pigott
Mark Clark	http://en.wikipedia.org/wiki/Mark_Wayne_Clark
Mark Consuelos	http://en.wikipedia.org/wiki/Mark_Consuelos
Mark Critz	http://en.wikipedia.org/wiki/Mark_Critz
Mark Cuban	http://en.wikipedia.org/wiki/Mark_Cuban
Mark D. Siljander	http://en.wikipedia.org/wiki/Mark_D._Siljander
Mark Dacascos	http://en.wikipedia.org/wiki/Mark_Dacascos
Mark David Chapman	http://en.wikipedia.org/wiki/Mark_David_Chapman
Mark Dayton	http://en.wikipedia.org/wiki/Mark_Dayton
Mark DeBarge	http://en.wikipedia.org/wiki/Mark_DeBarge
Mark Durkan	http://en.wikipedia.org/wiki/Mark_Durkan
Mark E. Smith	http://en.wikipedia.org/wiki/Mark_E._Smith
Mark Eitzel	http://en.wikipedia.org/wiki/Mark_Eitzel
Mark Feuerstein	http://en.wikipedia.org/wiki/Mark_Feuerstein
Mark Field	http://en.wikipedia.org/wiki/Mark_Field
Mark Foley	http://en.wikipedia.org/wiki/Mark_Foley
Mark Francois	http://en.wikipedia.org/wiki/Mark_Francois
Mark Fuhrman	http://en.wikipedia.org/wiki/Mark_Fuhrman
Mark Garnier	http://en.wikipedia.org/wiki/Mark_Garnier
Mark Gastineau	http://en.wikipedia.org/wiki/Mark_Gastineau
Mark Goddard	http://en.wikipedia.org/wiki/Mark_Goddard
Mark Green	http://en.wikipedia.org/wiki/Mark_Andrew_Green
Mark Haddon	http://en.wikipedia.org/wiki/Mark_Haddon
Mark Hamill	http://en.wikipedia.org/wiki/Mark_Hamill
Mark Harmon	http://en.wikipedia.org/wiki/Mark_Harmon
Mark Harper	http://en.wikipedia.org/wiki/Mark_Harper
Mark Hatfield	http://en.wikipedia.org/wiki/Mark_Hatfield
Mark Helprin	http://en.wikipedia.org/wiki/Mark_Helprin
Mark Hendrick	http://en.wikipedia.org/wiki/Mark_Hendrick
Mark Hoban	http://en.wikipedia.org/wiki/Mark_Hoban
Mark Hoppus	http://en.wikipedia.org/wiki/Mark_Hoppus
Mark Hunter	http://en.wikipedia.org/wiki/Mark_Hunter_(politician)
Mark Kennedy	http://en.wikipedia.org/wiki/Mark_Kennedy_(politician)
Mark Kirk	http://en.wikipedia.org/wiki/Mark_Kirk
Mark Knopfler	http://en.wikipedia.org/wiki/Mark_Knopfler
Mark Kozelek	http://en.wikipedia.org/wiki/Mark_Kozelek
Mark L. Lester	http://en.wikipedia.org/wiki/Mark_L._Lester
Mark Lancaster	http://en.wikipedia.org/wiki/Mark_Lancaster
Mark Lanegan	http://en.wikipedia.org/wiki/Mark_Lanegan
Mark Lazarowicz	http://en.wikipedia.org/wiki/Mark_Lazarowicz
Mark Lester	http://en.wikipedia.org/wiki/Mark_Lester
Mark Leyner	http://en.wikipedia.org/wiki/Mark_Leyner
Mark McGrath	http://en.wikipedia.org/wiki/Mark_McGrath
Mark McGwire	http://en.wikipedia.org/wiki/Mark_McGwire
Mark McKinney	http://en.wikipedia.org/wiki/Mark_McKinney
Mark Menzies	http://en.wikipedia.org/wiki/Mark_Menzies
Mark Millar	http://en.wikipedia.org/wiki/Mark_Millar
Mark Mothersbaugh	http://en.wikipedia.org/wiki/Mark_Mothersbaugh
Mark O. Hatfield	http://en.wikipedia.org/wiki/Mark_O._Hatfield
Mark Pauline	http://en.wikipedia.org/wiki/Mark_Pauline
Mark Pawsey	http://en.wikipedia.org/wiki/Mark_Pawsey
Mark Philippoussis	http://en.wikipedia.org/wiki/Mark_Philippoussis
Mark Prisk	http://en.wikipedia.org/wiki/Mark_Prisk
Mark Pritchard	http://en.wikipedia.org/wiki/Mark_Pritchard_(politician)
Mark Pryor	http://en.wikipedia.org/wiki/Mark_Pryor
Mark R. Hughes	http://en.wikipedia.org/wiki/Mark_R._Hughes
Mark Reckless	http://en.wikipedia.org/wiki/Mark_Reckless
Mark Roberts	http://en.wikipedia.org/wiki/Mark_Roberts_(streaker)
Mark Roberts	http://en.wikipedia.org/wiki/Mark_Roberts_%28footballer_born_1983%29
Mark Robson	http://en.wikipedia.org/wiki/Mark_Robson
Mark Roth	http://en.wikipedia.org/wiki/Mark_Roth
Mark Rothko	http://en.wikipedia.org/wiki/Mark_Rothko
Mark Ruffalo	http://en.wikipedia.org/wiki/Mark_Ruffalo
Mark Russell	http://en.wikipedia.org/wiki/Mark_Russell
Mark Rydell	http://en.wikipedia.org/wiki/Mark_Rydell
Mark S. Schweiker	http://en.wikipedia.org/wiki/Mark_S._Schweiker
Mark Sandrich	http://en.wikipedia.org/wiki/Mark_Sandrich
Mark Sanford	http://en.wikipedia.org/wiki/Mark_Sanford
Mark Sanford	http://en.wikipedia.org/wiki/Mark_Sanford
Mark Schauer	http://en.wikipedia.org/wiki/Mark_Schauer
Mark Shields	http://en.wikipedia.org/wiki/Mark_Shields
Mark Simmonds	http://en.wikipedia.org/wiki/Mark_Simmonds
Mark Souder	http://en.wikipedia.org/wiki/Mark_Souder
Mark Spencer	http://en.wikipedia.org/wiki/Mark_Spencer_(politician)
Mark Spitz	http://en.wikipedia.org/wiki/Mark_Spitz
Mark Strand	http://en.wikipedia.org/wiki/Mark_Strand
Mark Tami	http://en.wikipedia.org/wiki/Mark_Tami
Mark Tapio Kines	http://en.wikipedia.org/wiki/Mark_Tapio_Kines
Mark Thatcher	http://en.wikipedia.org/wiki/Mark_Thatcher
Mark Twain	http://en.wikipedia.org/wiki/Mark_Twain
Mark Udall	http://en.wikipedia.org/wiki/Mark_Udall
Mark Van Doren	http://en.wikipedia.org/wiki/Mark_Van_Doren
Mark Wahlberg	http://en.wikipedia.org/wiki/Mark_Wahlberg
Mark Warner	http://en.wikipedia.org/wiki/Mark_Warner
Mark Williams	http://en.wikipedia.org/wiki/Mark_Williams_(politician)
Mark Zuckerberg	http://en.wikipedia.org/wiki/Mark_Zuckerberg
Markie Post	http://en.wikipedia.org/wiki/Markie_Post
Mark-Paul Gosselaar	http://en.wikipedia.org/wiki/Mark-Paul_Gosselaar
Marla Gibbs	http://en.wikipedia.org/wiki/Marla_Gibbs
Marla Maples	http://en.wikipedia.org/wiki/Marla_Maples
Marla Sokoloff	http://en.wikipedia.org/wiki/Marla_Sokoloff
Marlee Matlin	http://en.wikipedia.org/wiki/Marlee_Matlin
Marlene Dietrich	http://en.wikipedia.org/wiki/Marlene_Dietrich
Marl�ne Jobert	http://en.wikipedia.org/wiki/Marl%E8ne_Jobert
Marlin Fitzwater	http://en.wikipedia.org/wiki/Marlin_Fitzwater
Marlin Perkins	http://en.wikipedia.org/wiki/Marlin_Perkins
Marlo Thomas	http://en.wikipedia.org/wiki/Marlo_Thomas
Marlon Brando	http://en.wikipedia.org/wiki/Marlon_Brando
Marlon Jackson	http://en.wikipedia.org/wiki/Marlon_Jackson
Marlon Wayans	http://en.wikipedia.org/wiki/Marlon_Wayans
Marques Houston	http://en.wikipedia.org/wiki/Marques_Houston
Marquis de Condorcet	http://en.wikipedia.org/wiki/Marquis_de_Condorcet
Marquis de Lafayette	http://en.wikipedia.org/wiki/Marquis_de_Lafayette
Marquis de Sade	http://en.wikipedia.org/wiki/Marquis_de_Sade
Marsha Blackburn	http://en.wikipedia.org/wiki/Marsha_Blackburn
Marsha Mason	http://en.wikipedia.org/wiki/Marsha_Mason
Marsha Singh	http://en.wikipedia.org/wiki/Marsha_Singh
Marshall Applewhite	http://en.wikipedia.org/wiki/Marshall_Applewhite
Marshall Hall	http://en.wikipedia.org/wiki/Marshall_Hall_(physiologist)
Marshall Holman	http://en.wikipedia.org/wiki/Marshall_Holman
Marshall McLuhan	http://en.wikipedia.org/wiki/Marshall_McLuhan
Marshall O. Larsen	http://en.wikipedia.org/wiki/Marshall_Larsen
Marshall Sylver	http://en.wikipedia.org/wiki/Marshall_Sylver
Marta Kauffman	http://en.wikipedia.org/wiki/Marta_Kauffman
Marta Kristen	http://en.wikipedia.org/wiki/Marta_Kristen
Martha Coolidge	http://en.wikipedia.org/wiki/Martha_Coolidge
Martha Graham	http://en.wikipedia.org/wiki/Martha_Graham
Martha Grimes	http://en.wikipedia.org/wiki/Martha_Grimes
Martha Moxley	http://en.wikipedia.org/wiki/Martha_Moxley
Martha Nussbaum	http://en.wikipedia.org/wiki/Martha_Nussbaum
Martha Plimpton	http://en.wikipedia.org/wiki/Martha_Plimpton
Martha Quinn	http://en.wikipedia.org/wiki/Martha_Quinn
Martha Raddatz	http://en.wikipedia.org/wiki/Martha_Raddatz
Martha Raye	http://en.wikipedia.org/wiki/Martha_Raye
Martha Reeves	http://en.wikipedia.org/wiki/Martha_Reeves
Martha Stewart	http://en.wikipedia.org/wiki/Martha_Stewart
Martha Washington	http://en.wikipedia.org/wiki/Martha_Washington
Martin Agronsky	http://en.wikipedia.org/wiki/Martin_Agronsky
Martin Amis	http://en.wikipedia.org/wiki/Martin_Amis
Martin Balsam	http://en.wikipedia.org/wiki/Martin_Balsam
Martin Bashir	http://en.wikipedia.org/wiki/Martin_Bashir
Martin Bormann	http://en.wikipedia.org/wiki/Martin_Bormann
Martin Boyd	http://en.wikipedia.org/wiki/Martin_Boyd
Martin Brest	http://en.wikipedia.org/wiki/Martin_Brest
Martin Bryant	http://en.wikipedia.org/wiki/Martin_Bryant
Martin Buber	http://en.wikipedia.org/wiki/Martin_Buber
Martin Bucer	http://en.wikipedia.org/wiki/Martin_Bucer
Martin Caton	http://en.wikipedia.org/wiki/Martin_Caton
Martin Chemnitz	http://en.wikipedia.org/wiki/Martin_Chemnitz
Martin Denny	http://en.wikipedia.org/wiki/Martin_Denny
Martin Donovan	http://en.wikipedia.org/wiki/Martin_Donovan
Martin Feldstein	http://en.wikipedia.org/wiki/Martin_Feldstein
Martin Flavin	http://en.wikipedia.org/wiki/Martin_Flavin
Martin Fleischmann	http://en.wikipedia.org/wiki/Martin_Fleischmann
Martin Freeman	http://en.wikipedia.org/wiki/Martin_Freeman
Martin Frost	http://en.wikipedia.org/wiki/Martin_Frost
Martin Frost	http://en.wikipedia.org/wiki/Martin_Frost
Martin Fry	http://en.wikipedia.org/wiki/Martin_Fry
Martin Garbus	http://en.wikipedia.org/wiki/Martin_Garbus
Martin Gardner	http://en.wikipedia.org/wiki/Martin_Gardner
Martin Gore	http://en.wikipedia.org/wiki/Martin_Gore
Martin Heidegger	http://en.wikipedia.org/wiki/Martin_Heidegger
Martin Heinrich	http://en.wikipedia.org/wiki/Martin_Heinrich
Martin Heinrich Klaproth	http://en.wikipedia.org/wiki/Martin_Heinrich_Klaproth
Martin Hellman	http://en.wikipedia.org/wiki/Martin_Hellman
Martin Henderson	http://en.wikipedia.org/wiki/Martin_Henderson
Martin Horwood	http://en.wikipedia.org/wiki/Martin_Horwood
Martin L. Perl	http://en.wikipedia.org/wiki/Martin_L._Perl
Martin Landau	http://en.wikipedia.org/wiki/Martin_Landau
Martin Lawrence	http://en.wikipedia.org/wiki/Martin_Lawrence
Martin Luther	http://en.wikipedia.org/wiki/Martin_Luther
Martin Luther King	http://en.wikipedia.org/wiki/Martin_Luther_King
Martin McGuinness	http://en.wikipedia.org/wiki/Martin_McGuinness
Martin Milner	http://en.wikipedia.org/wiki/Martin_Milner
Martin Mull	http://en.wikipedia.org/wiki/Martin_Mull
Martin Olav Sabo	http://en.wikipedia.org/wiki/Martin_Olav_Sabo
Martin O'Malley	http://en.wikipedia.org/wiki/Martin_O%27Malley
Martin O'Neill	http://en.wikipedia.org/wiki/Martin_O%27Neill
Martin Rev	http://en.wikipedia.org/wiki/Martin_Rev
Martin Ritt	http://en.wikipedia.org/wiki/Martin_Ritt
Martin Ryle	http://en.wikipedia.org/wiki/Martin_Ryle
Martin Sabo	http://en.wikipedia.org/wiki/Martin_Sabo
Martin Schmidt	http://en.wikipedia.org/wiki/Martin_Schmidt
Martin Schongauer	http://en.wikipedia.org/wiki/Martin_Schongauer
Martin Scorsese	http://en.wikipedia.org/wiki/Martin_Scorsese
Martin Sheen	http://en.wikipedia.org/wiki/Martin_Sheen
Martin Short	http://en.wikipedia.org/wiki/Martin_Short
Martin Shubik	http://en.wikipedia.org/wiki/Martin_Shubik
Mart�n Torrijos	http://en.wikipedia.org/wiki/Mart%EDn_Torrijos
Martin Tyler	http://en.wikipedia.org/wiki/Martin_Tyler
Martin Van Buren	http://en.wikipedia.org/wiki/Martin_Van_Buren
Martin Vickers	http://en.wikipedia.org/wiki/Martin_Vickers
Martin Waldseemuller	http://en.wikipedia.org/wiki/Martin_Waldseemuller
Martin Yan	http://en.wikipedia.org/wiki/Martin_Yan
Martina Hingis	http://en.wikipedia.org/wiki/Martina_Hingis
Martina McBride	http://en.wikipedia.org/wiki/Martina_McBride
Martina Navratilova	http://en.wikipedia.org/wiki/Martina_Navratilova
Martina Navratilova	http://en.wikipedia.org/wiki/Martina_Navratilova
Martine Dennis	http://en.wikipedia.org/wiki/Martine_Dennis
Martinus J.G. Veltman	http://en.wikipedia.org/wiki/Martinus_J.G._Veltman
Marty Allen	http://en.wikipedia.org/wiki/Marty_Allen_(comedian)
Marty Balin	http://en.wikipedia.org/wiki/Marty_Balin
Marty Feldman	http://en.wikipedia.org/wiki/Marty_Feldman
Marty Ingels	http://en.wikipedia.org/wiki/Marty_Ingels
Marty Krofft	http://en.wikipedia.org/wiki/Marty_Krofft
Marty Meehan	http://en.wikipedia.org/wiki/Marty_Meehan
Marty Robbins	http://en.wikipedia.org/wiki/Marty_Robbins
Marty Russo	http://en.wikipedia.org/wiki/Marty_Russo
Maruschka Detmers	http://en.wikipedia.org/wiki/Maruschka_Detmers
Marv Albert	http://en.wikipedia.org/wiki/Marv_Albert
Marv Wolfman	http://en.wikipedia.org/wiki/Marv_Wolfman
Marvin Bush	http://en.wikipedia.org/wiki/Marvin_Bush
Marvin Gaye	http://en.wikipedia.org/wiki/Marvin_Gaye
Marvin Hagler	http://en.wikipedia.org/wiki/Marvin_Hagler
Marvin Hamlisch	http://en.wikipedia.org/wiki/Marvin_Hamlisch
Marvin Harris	http://en.wikipedia.org/wiki/Marvin_Harris
Marvin Heemeyer	http://en.wikipedia.org/wiki/Marvin_Heemeyer
Marvin Kalb	http://en.wikipedia.org/wiki/Marvin_Kalb
Marvin Leath	http://en.wikipedia.org/wiki/Marvin_Leath
Marvin Minsky	http://en.wikipedia.org/wiki/Marvin_Minsky
Marvin Mitchelson	http://en.wikipedia.org/wiki/Marvin_Mitchelson
Marvin Olasky	http://en.wikipedia.org/wiki/Marvin_Olasky
Marvin Runyon	http://en.wikipedia.org/wiki/Marvin_Runyon
Mary Alden	http://en.wikipedia.org/wiki/Mary_Alden
Mary Ann Mobley	http://en.wikipedia.org/wiki/Mary_Ann_Mobley
Mary Antin	http://en.wikipedia.org/wiki/Mary_Antin
Mary Astor	http://en.wikipedia.org/wiki/Mary_Astor
Mary Austin	http://en.wikipedia.org/wiki/Mary_Austin
Mary Baker Eddy	http://en.wikipedia.org/wiki/Mary_Baker_Eddy
Mary Beth Hurt	http://en.wikipedia.org/wiki/Mary_Beth_Hurt
Mary Boland	http://en.wikipedia.org/wiki/Mary_Boland
Mary Bono	http://en.wikipedia.org/wiki/Mary_Bono
Mary Cassatt	http://en.wikipedia.org/wiki/Mary_Cassatt
Mary Chapin Carpenter	http://en.wikipedia.org/wiki/Mary_Chapin_Carpenter
Mary Cheney	http://en.wikipedia.org/wiki/Mary_Cheney
Mary Creagh	http://en.wikipedia.org/wiki/Mary_Creagh
Mary Crosby	http://en.wikipedia.org/wiki/Mary_Crosby
Mary Decker Slaney	http://en.wikipedia.org/wiki/Mary_Decker_Slaney
Mary Elizabeth Braddon	http://en.wikipedia.org/wiki/Mary_Elizabeth_Braddon
Mary Elizabeth Donaldson	http://en.wikipedia.org/wiki/Mary_Elizabeth_Donaldson
Mary Elizabeth Mastrantonio	http://en.wikipedia.org/wiki/Mary_Elizabeth_Mastrantonio
Mary Ellen Chase	http://en.wikipedia.org/wiki/Mary_Ellen_Chase
Mary Fallin	http://en.wikipedia.org/wiki/Mary_Fallin
Mary Flora Bell	http://en.wikipedia.org/wiki/Mary_Flora_Bell
Mary Frann	http://en.wikipedia.org/wiki/Mary_Frann
Mary Glindon	http://en.wikipedia.org/wiki/Mary_Glindon
Mary Hansen	http://en.wikipedia.org/wiki/Mary_Hansen
Mary Hart	http://en.wikipedia.org/wiki/Mary_Hart
Mary Higgins Clark	http://en.wikipedia.org/wiki/Mary_Higgins_Clark
Mary Hopkin	http://en.wikipedia.org/wiki/Mary_Hopkin
Mary I of Scotland	http://en.wikipedia.org/wiki/Mary_I_of_Scotland
Mary J. Blige	http://en.wikipedia.org/wiki/Mary_J._Blige
Mary Jo Kilroy	http://en.wikipedia.org/wiki/Mary_Jo_Kilroy
Mary Jo Kopechne	http://en.wikipedia.org/wiki/Mary_Jo_Kopechne
Mary Johnston	http://en.wikipedia.org/wiki/Mary_Johnston
Mary Karr	http://en.wikipedia.org/wiki/Mary_Karr
Mary Kay Letourneau	http://en.wikipedia.org/wiki/Mary_Kay_Letourneau
Mary Kay Place	http://en.wikipedia.org/wiki/Mary_Kay_Place
Mary Lambert	http://en.wikipedia.org/wiki/Mary_Lambert
Mary Landrieu	http://en.wikipedia.org/wiki/Mary_Landrieu
Mary Leakey	http://en.wikipedia.org/wiki/Mary_Leakey
Mary Lee Settle	http://en.wikipedia.org/wiki/Mary_Lee_Settle
Mary Lou Lord	http://en.wikipedia.org/wiki/Mary_Lou_Lord
Mary Lou Retton	http://en.wikipedia.org/wiki/Mary_Lou_Retton
Mary Lynn Rajskub	http://en.wikipedia.org/wiki/Mary_Lynn_Rajskub
Mary Lyon	http://en.wikipedia.org/wiki/Mary_Lyon
Mary MacLeod	http://en.wikipedia.org/wiki/Mary_MacLeod
Mary Magdalene	http://en.wikipedia.org/wiki/Mary_Magdalene
Mary Martin	http://en.wikipedia.org/wiki/Mary_Martin
Mary Matalin	http://en.wikipedia.org/wiki/Mary_Matalin
Mary McAleese	http://en.wikipedia.org/wiki/Mary_McAleese
Mary McCarthy	http://en.wikipedia.org/wiki/Mary_McCarthy_(author)
Mary McCormack	http://en.wikipedia.org/wiki/Mary_McCormack
Mary McDonnell	http://en.wikipedia.org/wiki/Mary_McDonnell
Mary McGrory	http://en.wikipedia.org/wiki/Mary_McGrory
Mary Midgley	http://en.wikipedia.org/wiki/Mary_Midgley
Mary Oliver	http://en.wikipedia.org/wiki/Mary_Oliver
Mary Pickford	http://en.wikipedia.org/wiki/Mary_Pickford
Mary Pierce	http://en.wikipedia.org/wiki/Mary_Pierce
Mary Renault	http://en.wikipedia.org/wiki/Mary_Renault
Mary Roberts Rinehart	http://en.wikipedia.org/wiki/Mary_Roberts_Rinehart
Mary Robinson	http://en.wikipedia.org/wiki/Mary_Robinson
Mary Rose Oakar	http://en.wikipedia.org/wiki/Mary_Rose_Oakar
Mary Rowlandson	http://en.wikipedia.org/wiki/Mary_Rowlandson
Mary Shelley	http://en.wikipedia.org/wiki/Mary_Shelley
Mary Steenburgen	http://en.wikipedia.org/wiki/Mary_Steenburgen
Mary Stuart Masterson	http://en.wikipedia.org/wiki/Mary_Stuart_Masterson
Mary Tamm	http://en.wikipedia.org/wiki/Mary_Tamm
Mary Timony	http://en.wikipedia.org/wiki/Mary_Timony
Mary Todd Lincoln	http://en.wikipedia.org/wiki/Mary_Todd_Lincoln
Mary Travers	http://en.wikipedia.org/wiki/Mary_Travers
Mary Tyler Moore	http://en.wikipedia.org/wiki/Mary_Tyler_Moore
Mary Wells	http://en.wikipedia.org/wiki/Mary_Wells
Mary Whitehouse	http://en.wikipedia.org/wiki/Mary_Whitehouse
Mary Wickes	http://en.wikipedia.org/wiki/Mary_Wickes
Mary Wilson	http://en.wikipedia.org/wiki/Mary_Wilson_(singer)
Mary Wollstonecraft	http://en.wikipedia.org/wiki/Mary_Wollstonecraft
Maryam d'Abo	http://en.wikipedia.org/wiki/Maryam_d%27Abo
Mary-Ellis Bunim	http://en.wikipedia.org/wiki/Mary-Ellis_Bunim
Mary-Kate Olsen	http://en.wikipedia.org/wiki/Mary-Kate_Olsen
Mary-Louise Parker	http://en.wikipedia.org/wiki/Mary-Louise_Parker
Masaharu Morimoto	http://en.wikipedia.org/wiki/Masaharu_Morimoto
Masahiko Kobe	http://en.wikipedia.org/wiki/Masahiko_Kobe
Masami Akita	http://en.wikipedia.org/wiki/Masami_Akita
Masamichi Amano	http://en.wikipedia.org/wiki/Masamichi_Amano
Masashi Amenomori	http://en.wikipedia.org/wiki/Masashi_Amenomori
Masatoshi Koshiba	http://en.wikipedia.org/wiki/Masatoshi_Koshiba
Mason Adams	http://en.wikipedia.org/wiki/Mason_Adams
Mason Locke Weems	http://en.wikipedia.org/wiki/Mason_Locke_Weems
Mason Reese	http://en.wikipedia.org/wiki/Mason_Reese
Masta Killa	http://en.wikipedia.org/wiki/Masta_Killa
Master P	http://en.wikipedia.org/wiki/Master_P
Masuo Amada	http://en.wikipedia.org/wiki/Masuo_Amada
Mata Hari	http://en.wikipedia.org/wiki/Mata_Hari
Mathew St. Patrick	http://en.wikipedia.org/wiki/Mathew_St._Patrick
Mathieu K�r�kou	http://en.wikipedia.org/wiki/Mathieu_K%E9r%E9kou
Matt Blunt	http://en.wikipedia.org/wiki/Matt_Blunt
Matt Blunt	http://en.wikipedia.org/wiki/Matt_Blunt
Matt Cameron	http://en.wikipedia.org/wiki/Matt_Cameron
Matt Craven	http://en.wikipedia.org/wiki/Matt_Craven
Matt Damon	http://en.wikipedia.org/wiki/Matt_Damon
Matt Dillon	http://en.wikipedia.org/wiki/Matt_Dillon
Matt Drudge	http://en.wikipedia.org/wiki/Matt_Drudge
Matt Frewer	http://en.wikipedia.org/wiki/Matt_Frewer
Matt Gonzalez	http://en.wikipedia.org/wiki/Matt_Gonzalez
Matt Groening	http://en.wikipedia.org/wiki/Matt_Groening
Matt Hale	http://en.wikipedia.org/wiki/Matthew_F._Hale
Matt Hasselbeck	http://en.wikipedia.org/wiki/Matt_Hasselbeck
Matt Lauer	http://en.wikipedia.org/wiki/Matt_Lauer
Matt LeBlanc	http://en.wikipedia.org/wiki/Matt_LeBlanc
Matt Letscher	http://en.wikipedia.org/wiki/Matt_Letscher
Matt Lucas	http://en.wikipedia.org/wiki/Matt_Lucas
Matt Salinger	http://en.wikipedia.org/wiki/Matt_Salinger
Matt Sharp	http://en.wikipedia.org/wiki/Matt_Sharp
Matt Sorum	http://en.wikipedia.org/wiki/Matt_Sorum
Matt Stone	http://en.wikipedia.org/wiki/Matt_Stone
Matteo Ricci	http://en.wikipedia.org/wiki/Matteo_Ricci
Matthew Arnold	http://en.wikipedia.org/wiki/Matthew_Arnold
Matthew Barney	http://en.wikipedia.org/wiki/Matthew_Barney
Matthew Bellamy	http://en.wikipedia.org/wiki/Matthew_Bellamy
Matthew Boulton	http://en.wikipedia.org/wiki/Matthew_Boulton
Matthew Bright	http://en.wikipedia.org/wiki/Matthew_Bright
Matthew Broderick	http://en.wikipedia.org/wiki/Matthew_Broderick
Matthew Cooper	http://en.wikipedia.org/wiki/Matthew_Cooper_(American_journalist)
Matthew Dowd	http://en.wikipedia.org/wiki/Matthew_Dowd
Matthew F. McHugh	http://en.wikipedia.org/wiki/Matthew_F._McHugh
Matthew Fox	http://en.wikipedia.org/wiki/Matthew_Fox_(actor)
Matthew Fox	http://en.wikipedia.org/wiki/Matthew_Fox_(priest)
Matthew G. Martinez	http://en.wikipedia.org/wiki/Matthew_G._Martinez
Matthew Goode	http://en.wikipedia.org/wiki/Matthew_Goode
Matthew Hancock	http://en.wikipedia.org/wiki/Matthew_Hancock
Matthew Henson	http://en.wikipedia.org/wiki/Matthew_Henson
Matthew Herbert	http://en.wikipedia.org/wiki/Matthew_Herbert
Matthew Holness	http://en.wikipedia.org/wiki/Matthew_Holness
Matthew J. Rinaldo	http://en.wikipedia.org/wiki/Matthew_J._Rinaldo
Matthew Josephson	http://en.wikipedia.org/wiki/Matthew_Josephson
Matthew K. Rose	http://en.wikipedia.org/wiki/Matthew_K._Rose
Matthew Laborteaux	http://en.wikipedia.org/wiki/Matthew_Laborteaux
Matthew Lawrence	http://en.wikipedia.org/wiki/Matthew_Lawrence
Matthew Lesko	http://en.wikipedia.org/wiki/Matthew_Lesko
Matthew Lillard	http://en.wikipedia.org/wiki/Matthew_Lillard
Matthew McConaughey	http://en.wikipedia.org/wiki/Matthew_McConaughey
Matthew McGrory	http://en.wikipedia.org/wiki/Matthew_McGrory
Matthew Miller	http://en.wikipedia.org/wiki/Matthew_Miller_(journalist)
Matthew Modine	http://en.wikipedia.org/wiki/Matthew_Modine
Matthew Offord	http://en.wikipedia.org/wiki/Matthew_Offord
Matthew Paris	http://en.wikipedia.org/wiki/Matthew_Paris
Matthew Parker	http://en.wikipedia.org/wiki/Matthew_Parker
Matthew Perry	http://en.wikipedia.org/wiki/Matthew_Perry
Matthew Perry	http://en.wikipedia.org/wiki/Matthew_C._Perry
Matthew Shepard	http://en.wikipedia.org/wiki/Matthew_Shepard
Matthew Shipp	http://en.wikipedia.org/wiki/Matthew_Shipp
Matthew Sweet	http://en.wikipedia.org/wiki/Matthew_Sweet
Matthew Vaughn	http://en.wikipedia.org/wiki/Matthew_Vaughn
Matthew Waterhouse	http://en.wikipedia.org/wiki/Matthew_Waterhouse
Matthew Webb	http://en.wikipedia.org/wiki/Matthew_Webb
Matthias Corvinus	http://en.wikipedia.org/wiki/Matthias_Corvinus
Matthias Gr�newald	http://en.wikipedia.org/wiki/Matthias_Gr%FCnewald
Matthias Sammer	http://en.wikipedia.org/wiki/Matthias_Sammer
Matti Nyk�nen	http://en.wikipedia.org/wiki/Matti_Nyk%E4nen
Matti Vanhanen	http://en.wikipedia.org/wiki/Matti_Vanhanen
Mattie Stepanek	http://en.wikipedia.org/wiki/Mattie_Stepanek
Maud Adams	http://en.wikipedia.org/wiki/Maud_Adams
Maumoon Abdul Gayoom	http://en.wikipedia.org/wiki/Maumoon_Abdul_Gayoom
Maura Tierney	http://en.wikipedia.org/wiki/Maura_Tierney
Maureen Dowd	http://en.wikipedia.org/wiki/Maureen_Dowd
Maureen Flannigan	http://en.wikipedia.org/wiki/Maureen_Flannigan
Maureen Lipman	http://en.wikipedia.org/wiki/Maureen_Lipman
Maureen McCormick	http://en.wikipedia.org/wiki/Maureen_McCormick
Maureen McGovern	http://en.wikipedia.org/wiki/Maureen_McGovern
Maureen O'Hara	http://en.wikipedia.org/wiki/Maureen_O%27Hara
Maureen O'Sullivan	http://en.wikipedia.org/wiki/Maureen_O%27Sullivan
Maureen Potter	http://en.wikipedia.org/wiki/Maureen_Potter
Maureen Reagan	http://en.wikipedia.org/wiki/Maureen_Reagan
Maureen Stapleton	http://en.wikipedia.org/wiki/Maureen_Stapleton
Maurice Benard	http://en.wikipedia.org/wiki/Maurice_Benard
Maurice Bishop	http://en.wikipedia.org/wiki/Maurice_Bishop
Maurice Chevalier	http://en.wikipedia.org/wiki/Maurice_Chevalier
Maurice Evans	http://en.wikipedia.org/wiki/Maurice_Evans_(actor)
Maurice Gibb	http://en.wikipedia.org/wiki/Maurice_Gibb
Maurice Hinchey	http://en.wikipedia.org/wiki/Maurice_Hinchey
Maurice Jarre	http://en.wikipedia.org/wiki/Maurice_Jarre
Maurice Leblanc	http://en.wikipedia.org/wiki/Maurice_Leblanc
Maurice Maeterlinck	http://en.wikipedia.org/wiki/Maurice_Maeterlinck
Maurice Merleau-Ponty	http://en.wikipedia.org/wiki/Maurice_Merleau-Ponty
Maurice of Nassau	http://en.wikipedia.org/wiki/Maurice_of_Nassau
Maurice of Saxony	http://en.wikipedia.org/wiki/Maurice_of_Saxony
Maurice Papon	http://en.wikipedia.org/wiki/Maurice_Papon
Maurice Prendergast	http://en.wikipedia.org/wiki/Maurice_Prendergast
Maurice R. Greenberg	http://en.wikipedia.org/wiki/Maurice_R._Greenberg
Maurice Ravel	http://en.wikipedia.org/wiki/Maurice_Ravel
Maurice Sendak	http://en.wikipedia.org/wiki/Maurice_Sendak
Maurice Wilkins	http://en.wikipedia.org/wiki/Maurice_Wilkins
Maurice, comte de Saxe	http://en.wikipedia.org/wiki/Maurice%2C_comte_de_Saxe
Mauricio Funes	http://en.wikipedia.org/wiki/Mauricio_Funes
Mauro Bolognini	http://en.wikipedia.org/wiki/Mauro_Bolognini
Maury Chaykin	http://en.wikipedia.org/wiki/Maury_Chaykin
Maury Povich	http://en.wikipedia.org/wiki/Maury_Povich
Mavis Gallant	http://en.wikipedia.org/wiki/Mavis_Gallant
Max Apple	http://en.wikipedia.org/wiki/Max_Apple
Max Baer	http://en.wikipedia.org/wiki/Max_Baer_(boxer)
Max Baer, Jr.	http://en.wikipedia.org/wiki/Max_Baer%2C_Jr.
Max Baucus	http://en.wikipedia.org/wiki/Max_Baucus
Max Baucus	http://en.wikipedia.org/wiki/Max_Baucus
Max Beerbohm	http://en.wikipedia.org/wiki/Max_Beerbohm
Max Born	http://en.wikipedia.org/wiki/Max_Born
Max Brod	http://en.wikipedia.org/wiki/Max_Brod
Max Bruch	http://en.wikipedia.org/wiki/Max_Bruch
Max Burns	http://en.wikipedia.org/wiki/Max_Burns
Max Cannon	http://en.wikipedia.org/wiki/Max_Cannon
Max Cavalera	http://en.wikipedia.org/wiki/Max_Cavalera
Max Cleland	http://en.wikipedia.org/wiki/Max_Cleland
Max Eastman	http://en.wikipedia.org/wiki/Max_Eastman
Max Ernst	http://en.wikipedia.org/wiki/Max_Ernst
Max F. Perutz	http://en.wikipedia.org/wiki/Max_F._Perutz
Max Frisch	http://en.wikipedia.org/wiki/Max_Frisch
Max Gail	http://en.wikipedia.org/wiki/Max_Gail
Max Geldray	http://en.wikipedia.org/wiki/Max_Geldray
Max Jacob	http://en.wikipedia.org/wiki/Max_Jacob
Max Lerner	http://en.wikipedia.org/wiki/Max_Lerner
Max Nordau	http://en.wikipedia.org/wiki/Max_Nordau
Max Perlich	http://en.wikipedia.org/wiki/Max_Perlich
Max Planck	http://en.wikipedia.org/wiki/Max_Planck
Max Roach	http://en.wikipedia.org/wiki/Max_Roach
Max Robinson	http://en.wikipedia.org/wiki/Max_Robinson
Max Sandlin	http://en.wikipedia.org/wiki/Max_Sandlin
Max Schmeling	http://en.wikipedia.org/wiki/Max_Schmeling
Max Stirner	http://en.wikipedia.org/wiki/Max_Stirner
Max van der Stoel	http://en.wikipedia.org/wiki/Max_van_der_Stoel
Max von Laue	http://en.wikipedia.org/wiki/Max_von_Laue
Max von Sydow	http://en.wikipedia.org/wiki/Max_von_Sydow
Max Weber	http://en.wikipedia.org/wiki/Max_Weber
Max Weinberg	http://en.wikipedia.org/wiki/Max_Weinberg
Max Wright	http://en.wikipedia.org/wiki/Max_Wright
Max Zorn	http://en.wikipedia.org/wiki/Max_Zorn
Maxfield Parrish	http://en.wikipedia.org/wiki/Maxfield_Parrish
Maxim Gorky	http://en.wikipedia.org/wiki/Maxim_Gorky
Maximilian I	http://en.wikipedia.org/wiki/Maximilian_I,_Holy_Roman_Emperor
Maximilian II	http://en.wikipedia.org/wiki/Maximilian_II,_Holy_Roman_Emperor
Maximilian Schell	http://en.wikipedia.org/wiki/Maximilian_Schell
Maximilian von Baden	http://en.wikipedia.org/wiki/Prince_Maximilian_of_Baden
Maximilien de B�thune	http://en.wikipedia.org/wiki/Maximilien_de_B%E9thune
Maxine Hong Kingston	http://en.wikipedia.org/wiki/Maxine_Hong_Kingston
Maxine Kumin	http://en.wikipedia.org/wiki/Maxine_Kumin
Maxine Waters	http://en.wikipedia.org/wiki/Maxine_Waters
Maxwell Anderson	http://en.wikipedia.org/wiki/Maxwell_Anderson
Maxwell Caulfield	http://en.wikipedia.org/wiki/Maxwell_Caulfield
May Miller	http://en.wikipedia.org/wiki/May_Miller
May Sarton	http://en.wikipedia.org/wiki/May_Sarton
May Swenson	http://en.wikipedia.org/wiki/May_Swenson
Maya Angelou	http://en.wikipedia.org/wiki/Maya_Angelou
Maya Lin	http://en.wikipedia.org/wiki/Maya_Lin
Maya Rudolph	http://en.wikipedia.org/wiki/Maya_Rudolph
Mayim Bialik	http://en.wikipedia.org/wiki/Mayim_Bialik
Maynard James Keenan	http://en.wikipedia.org/wiki/Maynard_James_Keenan
Mayo A. Shattuck III	http://en.wikipedia.org/wiki/Mayo_A._Shattuck_III
Mayo Thompson	http://en.wikipedia.org/wiki/Mayo_Thompson
Mazie Hirono	http://en.wikipedia.org/wiki/Mazie_Hirono
MC 900 Ft. Jesus	http://en.wikipedia.org/wiki/MC_900_Ft._Jesus
mc chris	http://en.wikipedia.org/wiki/mc_chris
MC Hammer	http://en.wikipedia.org/wiki/MC_Hammer
MC Lyte	http://en.wikipedia.org/wiki/MC_Lyte
MC Ren	http://en.wikipedia.org/wiki/MC_Ren
MC Serch	http://en.wikipedia.org/wiki/MC_Serch
McLean Stevenson	http://en.wikipedia.org/wiki/McLean_Stevenson
Meadowlark Lemon	http://en.wikipedia.org/wiki/Meadowlark_Lemon
Meagan Good	http://en.wikipedia.org/wiki/Meagan_Good
Meat Loaf	http://en.wikipedia.org/wiki/Meat_Loaf
Medgar Evers	http://en.wikipedia.org/wiki/Medgar_Evers
Meg Cabot	http://en.wikipedia.org/wiki/Meg_Cabot
Meg Foster	http://en.wikipedia.org/wiki/Meg_Foster
Meg Greenfield	http://en.wikipedia.org/wiki/Meg_Greenfield
Meg Hillier	http://en.wikipedia.org/wiki/Meg_Hillier
Meg Munn	http://en.wikipedia.org/wiki/Meg_Munn
Meg Ryan	http://en.wikipedia.org/wiki/Meg_Ryan
Meg Tilly	http://en.wikipedia.org/wiki/Meg_Tilly
Meg White	http://en.wikipedia.org/wiki/Meg_White
Meg Whitman	http://en.wikipedia.org/wiki/Meg_Whitman
Megan Follows	http://en.wikipedia.org/wiki/Megan_Follows
Megan Gallagher	http://en.wikipedia.org/wiki/Megan_Gallagher
Megan McCafferty	http://en.wikipedia.org/wiki/Megan_McCafferty
Megan Mullally	http://en.wikipedia.org/wiki/Megan_Mullally
Megawati Sukarnoputri	http://en.wikipedia.org/wiki/Megawati_Sukarnoputri
Mehmed I	http://en.wikipedia.org/wiki/Mehmed_I
Mehmed the Conqueror	http://en.wikipedia.org/wiki/Mehmed_the_Conqueror
Mehmet Ali Agca	http://en.wikipedia.org/wiki/Mehmet_Ali_Agca
Mehmet Ali Talat	http://en.wikipedia.org/wiki/Mehmet_Ali_Talat
Meindert Hobbema	http://en.wikipedia.org/wiki/Meindert_Hobbema
Meir Kahane	http://en.wikipedia.org/wiki/Meir_Kahane
Meister Eckhart	http://en.wikipedia.org/wiki/Meister_Eckhart
Mekhi Phifer	http://en.wikipedia.org/wiki/Mekhi_Phifer
Mel Blanc	http://en.wikipedia.org/wiki/Mel_Blanc
Mel Brooks	http://en.wikipedia.org/wiki/Mel_Brooks
Mel Carnahan	http://en.wikipedia.org/wiki/Mel_Carnahan
Mel Carter	http://en.wikipedia.org/wiki/Mel_Carter
Mel Collins	http://en.wikipedia.org/wiki/Mel_Collins
Mel Ferrer	http://en.wikipedia.org/wiki/Mel_Ferrer
Mel Gibson	http://en.wikipedia.org/wiki/Mel_Gibson
Mel Harris	http://en.wikipedia.org/wiki/Mel_Harris
Mel Karmazin	http://en.wikipedia.org/wiki/Mel_Karmazin
Mel Levine	http://en.wikipedia.org/wiki/Mel_Levine
Mel Martinez	http://en.wikipedia.org/wiki/Mel_Martinez
Mel Ott	http://en.wikipedia.org/wiki/Mel_Ott
Mel Reynolds	http://en.wikipedia.org/wiki/Mel_Reynolds
Mel Smith	http://en.wikipedia.org/wiki/Mel_Smith
Mel Stride	http://en.wikipedia.org/wiki/Mel_Stride
Mel Tillis	http://en.wikipedia.org/wiki/Mel_Tillis
Mel Torm�	http://en.wikipedia.org/wiki/Mel_Torm%E9
Mel Watt	http://en.wikipedia.org/wiki/Mel_Watt
Melanie B	http://en.wikipedia.org/wiki/Melanie_B
Melanie Blatt	http://en.wikipedia.org/wiki/Melanie_Blatt
Melanie C	http://en.wikipedia.org/wiki/Melanie_C
Melanie Chartoff	http://en.wikipedia.org/wiki/Melanie_Chartoff
Melanie Griffith	http://en.wikipedia.org/wiki/Melanie_Griffith
Melanie Lynskey	http://en.wikipedia.org/wiki/Melanie_Lynskey
Melanie Morgan	http://en.wikipedia.org/wiki/Melanie_Morgan
Melba Moore	http://en.wikipedia.org/wiki/Melba_Moore
Melchior Hofmann	http://en.wikipedia.org/wiki/Melchior_Hofmann
Melchiorre Gioja	http://en.wikipedia.org/wiki/Melchiorre_Gioja
Meles Zenawi	http://en.wikipedia.org/wiki/Meles_Zenawi
Melina Mercouri	http://en.wikipedia.org/wiki/Melina_Mercouri
Melinda Clarke	http://en.wikipedia.org/wiki/Melinda_Clarke
Melinda Gates	http://en.wikipedia.org/wiki/Melinda_Gates
Melissa Auf der Maur	http://en.wikipedia.org/wiki/Melissa_Auf_der_Maur
Melissa Bean	http://en.wikipedia.org/wiki/Melissa_Bean
Melissa Etheridge	http://en.wikipedia.org/wiki/Melissa_Etheridge
Melissa George	http://en.wikipedia.org/wiki/Melissa_George
Melissa Gilbert	http://en.wikipedia.org/wiki/Melissa_Gilbert
Melissa Hart	http://en.wikipedia.org/wiki/Melissa_Hart
Melissa Joan Hart	http://en.wikipedia.org/wiki/Melissa_Joan_Hart
Melissa Leo	http://en.wikipedia.org/wiki/Melissa_Leo
Melissa Manchester	http://en.wikipedia.org/wiki/Melissa_Manchester
Melissa Rivers	http://en.wikipedia.org/wiki/Melissa_Rivers
Melissa Sue Anderson	http://en.wikipedia.org/wiki/Melissa_Sue_Anderson
Melody Patterson	http://en.wikipedia.org/wiki/Melody_Patterson
Melvil Dewey	http://en.wikipedia.org/wiki/Melvil_Dewey
Melvin Belli	http://en.wikipedia.org/wiki/Melvin_Belli
Melvin Calvin	http://en.wikipedia.org/wiki/Melvin_Calvin
Melvin Franklin	http://en.wikipedia.org/wiki/Melvin_Franklin
Melvin J. Lasky	http://en.wikipedia.org/wiki/Melvin_J._Lasky
Melvin Laird	http://en.wikipedia.org/wiki/Melvin_Laird
Melvin Price	http://en.wikipedia.org/wiki/Melvin_Price
Melvin Schwartz	http://en.wikipedia.org/wiki/Melvin_Schwartz
Melvin Van Peebles	http://en.wikipedia.org/wiki/Melvin_Van_Peebles
Melvyn Bragg	http://en.wikipedia.org/wiki/Melvyn_Bragg
Melvyn Douglas	http://en.wikipedia.org/wiki/Melvyn_Douglas
Melyssa Ade	http://en.wikipedia.org/wiki/Melyssa_Ade
Memphis Bleek	http://en.wikipedia.org/wiki/Memphis_Bleek
Mena Suvari	http://en.wikipedia.org/wiki/Mena_Suvari
Menachem Begin	http://en.wikipedia.org/wiki/Menachem_Begin
Menasseh ben Israel	http://en.wikipedia.org/wiki/Menasseh_ben_Israel
Menno Simons	http://en.wikipedia.org/wiki/Menno_Simons
Menzies Campbell	http://en.wikipedia.org/wiki/Menzies_Campbell
Mercedes Lackey	http://en.wikipedia.org/wiki/Mercedes_Lackey
Mercedes McCambridge	http://en.wikipedia.org/wiki/Mercedes_McCambridge
Mercedes Ruehl	http://en.wikipedia.org/wiki/Mercedes_Ruehl
Mercer Reynolds	http://en.wikipedia.org/wiki/Mercer_Reynolds
Mercy Otis Warren	http://en.wikipedia.org/wiki/Mercy_Otis_Warren
Meredith Baxter	http://en.wikipedia.org/wiki/Meredith_Baxter
Meredith MacRae	http://en.wikipedia.org/wiki/Meredith_MacRae
Meredith Monk	http://en.wikipedia.org/wiki/Meredith_Monk
Meredith Monroe	http://en.wikipedia.org/wiki/Meredith_Monroe
Meredith Vieira	http://en.wikipedia.org/wiki/Meredith_Vieira
Merhan Karimi Nasseri	http://en.wikipedia.org/wiki/Merhan_Karimi_Nasseri
Meridel Le Sueur	http://en.wikipedia.org/wiki/Meridel_Le_Sueur
Meriwether Lewis	http://en.wikipedia.org/wiki/Meriwether_Lewis
Merl Saunders	http://en.wikipedia.org/wiki/Merl_Saunders
Merle Haggard	http://en.wikipedia.org/wiki/Merle_Haggard
Merle Oberon	http://en.wikipedia.org/wiki/Merle_Oberon
Merle Travis	http://en.wikipedia.org/wiki/Merle_Travis
Merlin Olsen	http://en.wikipedia.org/wiki/Merlin_Olsen
Merlin Santana	http://en.wikipedia.org/wiki/Merlin_Santana
Merrie Spaeth	http://en.wikipedia.org/wiki/Merrie_Spaeth
Merry Anders	http://en.wikipedia.org/wiki/Merry_Anders
Merv Griffin	http://en.wikipedia.org/wiki/Merv_Griffin
Mervat Amin	http://en.wikipedia.org/wiki/Mervat_Amin
Mervyn LeRoy	http://en.wikipedia.org/wiki/Mervyn_LeRoy
Mervyn M. Dymally	http://en.wikipedia.org/wiki/Mervyn_M._Dymally
Mervyn Peake	http://en.wikipedia.org/wiki/Mervyn_Peake
Meryl Streep	http://en.wikipedia.org/wiki/Meryl_Streep
Me'Shell Ndeg�Ocello	http://en.wikipedia.org/wiki/Me%27Shell_Ndeg%E9Ocello
Method Man	http://en.wikipedia.org/wiki/Method_Man
Meyer Lansky	http://en.wikipedia.org/wiki/Meyer_Lansky
Meyer Levin	http://en.wikipedia.org/wiki/Meyer_Levin
MF Doom	http://en.wikipedia.org/wiki/MF_Doom
MH Abrams	http://en.wikipedia.org/wiki/MH_Abrams
Mia Farrow	http://en.wikipedia.org/wiki/Mia_Farrow
Mia Hamm	http://en.wikipedia.org/wiki/Mia_Hamm
Mia Kirshner	http://en.wikipedia.org/wiki/Mia_Kirshner
Mia Sara	http://en.wikipedia.org/wiki/Mia_Sara
Mia Tyler	http://en.wikipedia.org/wiki/Mia_Tyler
Mic Geronimo	http://en.wikipedia.org/wiki/Mic_Geronimo
Michael A. Andrews	http://en.wikipedia.org/wiki/Michael_A._Andrews
Michael Addis	http://en.wikipedia.org/wiki/Michael_Addis
Michael Allinson	http://en.wikipedia.org/wiki/Michael_Allinson
Michael Anderson	http://en.wikipedia.org/wiki/Michael_Anderson_(director)
Michael Andretti	http://en.wikipedia.org/wiki/Michael_Andretti
Michael Angarano	http://en.wikipedia.org/wiki/Michael_Angarano
Michael Ansara	http://en.wikipedia.org/wiki/Michael_Ansara
Michael Anthony	http://en.wikipedia.org/wiki/Michael_Anthony_(musician)
Michael Anthony	http://en.wikipedia.org/wiki/Michael_Anthony_(author)
Michael Apted	http://en.wikipedia.org/wiki/Michael_Apted
Michael Arcuri	http://en.wikipedia.org/wiki/Michael_Arcuri
Michael Aspel	http://en.wikipedia.org/wiki/Michael_Aspel
Michael Badalucco	http://en.wikipedia.org/wiki/Michael_Badalucco
Michael Baius	http://en.wikipedia.org/wiki/Michael_Baius
Michael Bay	http://en.wikipedia.org/wiki/Michael_Bay
Michael Behe	http://en.wikipedia.org/wiki/Michael_Behe
Michael Bennet	http://en.wikipedia.org/wiki/Michael_Bennet
Michael Bergin	http://en.wikipedia.org/wiki/Michael_Bergin
Michael Berryman	http://en.wikipedia.org/wiki/Michael_Berryman
Michael Beschloss	http://en.wikipedia.org/wiki/Michael_Beschloss
Michael Biehn	http://en.wikipedia.org/wiki/Michael_Biehn
Michael Bilirakis	http://en.wikipedia.org/wiki/Michael_Bilirakis
Michael Bilirakis	http://en.wikipedia.org/wiki/Michael_Bilirakis
Michael Bloomberg	http://en.wikipedia.org/wiki/Michael_Bloomberg
Michael Boatman	http://en.wikipedia.org/wiki/Michael_Boatman
Michael Bolton	http://en.wikipedia.org/wiki/Michael_Bolton
Michael Bubl�	http://en.wikipedia.org/wiki/Michael_Bubl%E9
Michael Burgess	http://en.wikipedia.org/wiki/Michael_C._Burgess
Michael C. Hall	http://en.wikipedia.org/wiki/Michael_C._Hall
Michael C. Williams	http://en.wikipedia.org/wiki/Michael_C._Williams
Michael Caine	http://en.wikipedia.org/wiki/Michael_Caine
Michael Carroll	http://en.wikipedia.org/wiki/Michael_Carroll_(lottery_winner)
Michael Cera	http://en.wikipedia.org/wiki/Michael_Cera
Michael Chabon	http://en.wikipedia.org/wiki/Michael_Chabon
Michael Chapman	http://en.wikipedia.org/wiki/Michael_Chapman_(musician)
Michael Chertoff	http://en.wikipedia.org/wiki/Michael_Chertoff
Michael Chiklis	http://en.wikipedia.org/wiki/Michael_Chiklis
Michael Chow Man-Kin	http://en.wikipedia.org/wiki/Michael_Chow_Man-Kin
Michael Cimino	http://en.wikipedia.org/wiki/Michael_Cimino
Michael Clarke Duncan	http://en.wikipedia.org/wiki/Michael_Clarke_Duncan
Michael Collins	http://en.wikipedia.org/wiki/Michael_Collins_(astronaut)
Michael Collins	http://en.wikipedia.org/wiki/Michael_Collins_(Irish_leader)
Michael Connarty	http://en.wikipedia.org/wiki/Michael_Connarty
Michael Copps	http://en.wikipedia.org/wiki/Michael_Copps
Michael Crapo	http://en.wikipedia.org/wiki/Michael_Crapo
Michael Crawford	http://en.wikipedia.org/wiki/Michael_Crawford
Michael Crichton	http://en.wikipedia.org/wiki/Michael_Crichton
Michael Cunningham	http://en.wikipedia.org/wiki/Michael_Cunningham
Michael Curtiz	http://en.wikipedia.org/wiki/Michael_Curtiz
Michael D. Barnes	http://en.wikipedia.org/wiki/Michael_D._Barnes
Michael D. Brown	http://en.wikipedia.org/wiki/Michael_D._Brown
Michael Davitt	http://en.wikipedia.org/wiki/Michael_Davitt
Michael Deaver	http://en.wikipedia.org/wiki/Michael_Deaver
Michael DeBakey	http://en.wikipedia.org/wiki/Michael_DeBakey
Michael Dell	http://en.wikipedia.org/wiki/Michael_Dell
Michael DeLorenzo	http://en.wikipedia.org/wiki/Michael_DeLorenzo
Michael Dorn	http://en.wikipedia.org/wiki/Michael_Dorn
Michael Douglas	http://en.wikipedia.org/wiki/Michael_Douglas
Michael Drosnin	http://en.wikipedia.org/wiki/Michael_Drosnin
Michael Dugher	http://en.wikipedia.org/wiki/Michael_Dugher
Michael Dukakis	http://en.wikipedia.org/wiki/Michael_Dukakis
Michael E. Brown	http://en.wikipedia.org/wiki/Michael_E._Brown
Michael E. Capuano	http://en.wikipedia.org/wiki/Michael_E._Capuano
Michael Ealy	http://en.wikipedia.org/wiki/Michael_Ealy
Michael Easley	http://en.wikipedia.org/wiki/Mike_Easley
Michael Eisner	http://en.wikipedia.org/wiki/Michael_Eisner
Michael Ellis	http://en.wikipedia.org/wiki/Michael_Ellis_(British_politician)
Michael Enzi	http://en.wikipedia.org/wiki/Michael_Enzi
Michael Fabricant	http://en.wikipedia.org/wiki/Michael_Fabricant
Michael Fallon	http://en.wikipedia.org/wiki/Michael_Fallon
Michael Faraday	http://en.wikipedia.org/wiki/Michael_Faraday
Michael Feinstein	http://en.wikipedia.org/wiki/Michael_Feinstein
Michael Ferguson	http://en.wikipedia.org/wiki/Mike_Ferguson_(New_Jersey_politician)
Michael Fishman	http://en.wikipedia.org/wiki/Michael_Fishman
Michael Flatley	http://en.wikipedia.org/wiki/Michael_Flatley
Michael Franti	http://en.wikipedia.org/wiki/Michael_Franti
Michael G. Morris	http://en.wikipedia.org/wiki/Michael_G._Morris
Michael G. Mullen	http://en.wikipedia.org/wiki/Michael_G._Mullen
Michael G. Oxley	http://en.wikipedia.org/wiki/Michael_G._Oxley
Michael Gambon	http://en.wikipedia.org/wiki/Michael_Gambon
Michael Gerson	http://en.wikipedia.org/wiki/Michael_Gerson
Michael Giles	http://en.wikipedia.org/wiki/Michael_Giles
Michael Gira	http://en.wikipedia.org/wiki/Michael_Gira
Michael Gough	http://en.wikipedia.org/wiki/Michael_Gough
Michael Gove	http://en.wikipedia.org/wiki/Michael_Gove
Michael Gross	http://en.wikipedia.org/wiki/Michael_Gross_(actor)
Michael H. Jordan	http://en.wikipedia.org/wiki/Michael_H._Jordan
Michael Harrington	http://en.wikipedia.org/wiki/Michael_Harrington
Michael Haydn	http://en.wikipedia.org/wiki/Michael_Haydn
Michael Hoffman	http://en.wikipedia.org/wiki/Michael_Hoffman_(American_director)
Michael Hordern	http://en.wikipedia.org/wiki/Michael_Hordern
Michael Howard	http://en.wikipedia.org/wiki/Michael_Howard
Michael Huffington	http://en.wikipedia.org/wiki/Michael_Huffington
Michael Hutchence	http://en.wikipedia.org/wiki/Michael_Hutchence
Michael I. Sovern	http://en.wikipedia.org/wiki/Michael_I._Sovern
Michael Ian Black	http://en.wikipedia.org/wiki/Michael_Ian_Black
Michael Ignatieff	http://en.wikipedia.org/wiki/Michael_Ignatieff
Michael Imperioli	http://en.wikipedia.org/wiki/Michael_Imperioli
Michael Ironside	http://en.wikipedia.org/wiki/Michael_Ironside
Michael Irvin	http://en.wikipedia.org/wiki/Michael_Irvin
Michael Isikoff	http://en.wikipedia.org/wiki/Michael_Isikoff
Michael Ivins	http://en.wikipedia.org/wiki/Michael_Ivins
Michael J. Fox	http://en.wikipedia.org/wiki/Michael_J._Fox
Michael J. Jackson	http://en.wikipedia.org/wiki/Mike_Jackson_(auto)
Michael J. Nelson	http://en.wikipedia.org/wiki/Michael_J._Nelson
Michael Jackson	http://en.wikipedia.org/wiki/Michael_Jackson
Michael Jeffery	http://en.wikipedia.org/wiki/Michael_Jeffery
Michael Jeter	http://en.wikipedia.org/wiki/Michael_Jeter
Michael Johns	http://en.wikipedia.org/wiki/Michael_Johns_(executive)
Michael Jordan	http://en.wikipedia.org/wiki/Michael_Jordan
Michael Kearns	http://en.wikipedia.org/wiki/Michael_Kearns
Michael Keaton	http://en.wikipedia.org/wiki/Michael_Keaton
Michael Kelly	http://en.wikipedia.org/wiki/Michael_Kelly_(American_actor)
Michael Kidd	http://en.wikipedia.org/wiki/Michael_Kidd
Michael Kinsley	http://en.wikipedia.org/wiki/Michael_Kinsley
Michael Korda	http://en.wikipedia.org/wiki/Michael_Korda
Michael L. Eskew	http://en.wikipedia.org/wiki/Michael_L._Eskew
Michael L. Strang	http://en.wikipedia.org/wiki/Michael_L._Strang
Michael Landon	http://en.wikipedia.org/wiki/Michael_Landon
Michael Learned	http://en.wikipedia.org/wiki/Michael_Learned
Michael Ledeen	http://en.wikipedia.org/wiki/Michael_Ledeen
Michael Lewis	http://en.wikipedia.org/wiki/Michael_Lewis_(author)
Michael Madsen	http://en.wikipedia.org/wiki/Michael_Madsen
Michael Mann	http://en.wikipedia.org/wiki/Michael_Mann_(director)
Michael Mantler	http://en.wikipedia.org/wiki/Michael_Mantler
Michael Markowitz	http://en.wikipedia.org/wiki/Michael_Markowitz
Michael McCann	http://en.wikipedia.org/wiki/Michael_McCann_(politician)
Michael McCaul	http://en.wikipedia.org/wiki/Michael_McCaul
Michael McClure	http://en.wikipedia.org/wiki/Michael_McClure
Michael McDermott	http://en.wikipedia.org/wiki/Wakefield_Massacre
Michael McDonald	http://en.wikipedia.org/wiki/Michael_McDonald_(actor)
Michael McDonald	http://en.wikipedia.org/wiki/Michael_McDonald_(singer)
Michael McKean	http://en.wikipedia.org/wiki/Michael_McKean
Michael McMahon	http://en.wikipedia.org/wiki/Michael_McMahon
Michael McNulty	http://en.wikipedia.org/wiki/Michael_McNulty
Michael Meacher	http://en.wikipedia.org/wiki/Michael_Meacher
Michael Medved	http://en.wikipedia.org/wiki/Michael_Medved
Michael Melvill	http://en.wikipedia.org/wiki/Michael_Melvill
Michael Michaud	http://en.wikipedia.org/wiki/Michael_Michaud
Michael Michele	http://en.wikipedia.org/wiki/Michael_Michele
Michael Milken	http://en.wikipedia.org/wiki/Michael_Milken
Michael Moorcock	http://en.wikipedia.org/wiki/Michael_Moorcock
Michael Moore	http://en.wikipedia.org/wiki/Michael_Moore
Michael Moore	http://en.wikipedia.org/wiki/Michael_Moore_(UK_politician)
Michael Moriarty	http://en.wikipedia.org/wiki/Michael_Moriarty
Michael Murphy	http://en.wikipedia.org/wiki/Michael_Murphy_(actor)
Michael Musto	http://en.wikipedia.org/wiki/Michael_Musto
Michael Newdow	http://en.wikipedia.org/wiki/Michael_Newdow
Michael Ninn	http://en.wikipedia.org/wiki/Michael_Ninn
Michael Nouri	http://en.wikipedia.org/wiki/Michael_Nouri
Michael Novak	http://en.wikipedia.org/wiki/Michael_Novak
Michael O. Leavitt	http://en.wikipedia.org/wiki/Michael_O._Leavitt
Michael O'Keefe	http://en.wikipedia.org/wiki/Michael_O%27Keefe
Michael Ondaatje	http://en.wikipedia.org/wiki/Michael_Ondaatje
Michael Ontkean	http://en.wikipedia.org/wiki/Michael_Ontkean
Michael Ovitz	http://en.wikipedia.org/wiki/Michael_Ovitz
Michael Owen	http://en.wikipedia.org/wiki/Michael_Owen
Michael Oxley	http://en.wikipedia.org/wiki/Michael_Oxley
Michael Palin	http://en.wikipedia.org/wiki/Michael_Palin
Michael Par�	http://en.wikipedia.org/wiki/Michael_Par%E9
Michael Parks	http://en.wikipedia.org/wiki/Michael_Parks
Michael Patrick Jann	http://en.wikipedia.org/wiki/Michael_Patrick_Jann
Michael Paul Chan	http://en.wikipedia.org/wiki/Michael_Paul_Chan
Michael Penn	http://en.wikipedia.org/wiki/Michael_Penn
Michael Peterson	http://en.wikipedia.org/wiki/Michael_Peterson_(author)
Michael Phelps	http://en.wikipedia.org/wiki/Michael_Phelps
Michael Pitt	http://en.wikipedia.org/wiki/Michael_Pitt
Michael Porter	http://en.wikipedia.org/wiki/Michael_Porter
Michael Portillo	http://en.wikipedia.org/wiki/Michael_Portillo
Michael Powell	http://en.wikipedia.org/wiki/Michael_Powell_(politician)
Michael Powell	http://en.wikipedia.org/wiki/Michael_Powell_(director)
Michael Quigley	http://en.wikipedia.org/wiki/Michael_Quigley
Michael Rapaport	http://en.wikipedia.org/wiki/Michael_Rapaport
Michael Reagan	http://en.wikipedia.org/wiki/Michael_Reagan
Michael Redgrave	http://en.wikipedia.org/wiki/Michael_Redgrave
Michael Rennie	http://en.wikipedia.org/wiki/Michael_Rennie
Michael Richards	http://en.wikipedia.org/wiki/Michael_Richards
Michael Ritchie	http://en.wikipedia.org/wiki/Michael_Ritchie_(film_director)
Michael Rosenbaum	http://en.wikipedia.org/wiki/Michael_Rosenbaum
Michael Rumaker	http://en.wikipedia.org/wiki/Michael_Rumaker
Michael S. Steele	http://en.wikipedia.org/wiki/Michael_S._Steele
Michael Sandison	http://en.wikipedia.org/wiki/Michael_Sandison
Michael Sarrazin	http://en.wikipedia.org/wiki/Michael_Sarrazin
Michael Savage	http://en.wikipedia.org/wiki/Michael_Savage_(commentator)
Michael Schenker	http://en.wikipedia.org/wiki/Michael_Schenker
Michael Scheuer	http://en.wikipedia.org/wiki/Michael_Scheuer
Michael Schiavo	http://en.wikipedia.org/wiki/Michael_Schiavo
Michael Schumacher	http://en.wikipedia.org/wiki/Michael_Schumacher
Michael Servetus	http://en.wikipedia.org/wiki/Michael_Servetus
Michael Shaara	http://en.wikipedia.org/wiki/Michael_Shaara
Michael Shanks	http://en.wikipedia.org/wiki/Michael_Shanks
Michael Sheen	http://en.wikipedia.org/wiki/Michael_Sheen
Michael Shermer	http://en.wikipedia.org/wiki/Michael_Shermer
Michael Showalter	http://en.wikipedia.org/wiki/Michael_Showalter
Michael Skakel	http://en.wikipedia.org/wiki/Michael_Skakel
Michael Smith	http://en.wikipedia.org/wiki/Michael_Smith_(chemist)
Michael Spindler	http://en.wikipedia.org/wiki/Michael_Spindler
Michael Spinks	http://en.wikipedia.org/wiki/Michael_Spinks
Michael Starr	http://en.wikipedia.org/wiki/Michael_Starr
Michael Steele	http://en.wikipedia.org/wiki/Michael_Steele_(musician)
Michael Stipe	http://en.wikipedia.org/wiki/Michael_Stipe
Michael Storm	http://en.wikipedia.org/wiki/Michael_Storm
Michael T. Weiss	http://en.wikipedia.org/wiki/Michael_T._Weiss
Michael Turner	http://en.wikipedia.org/wiki/Mike_Turner
Michael V. Hayden	http://en.wikipedia.org/wiki/Michael_V._Hayden
Michael Vale	http://en.wikipedia.org/wiki/Michael_Vale
Michael Vartan	http://en.wikipedia.org/wiki/Michael_Vartan
Michael Vick	http://en.wikipedia.org/wiki/Michael_Vick
Michael Walzer	http://en.wikipedia.org/wiki/Michael_Walzer
Michael Warner	http://en.wikipedia.org/wiki/Michael_Warner
Michael Weatherly	http://en.wikipedia.org/wiki/Michael_Weatherly
Michael Welch	http://en.wikipedia.org/wiki/Michael_Welch_(actor)
Michael Wigglesworth	http://en.wikipedia.org/wiki/Michael_Wigglesworth
Michael Wilbon	http://en.wikipedia.org/wiki/Michael_Wilbon
Michael Wilding	http://en.wikipedia.org/wiki/Michael_Wilding_(actor)
Michael Williams	http://en.wikipedia.org/wiki/Michael_Williams_(actor)
Michael Wincott	http://en.wikipedia.org/wiki/Michael_Wincott
Michael Winner	http://en.wikipedia.org/wiki/Michael_Winner
Michael Winslow	http://en.wikipedia.org/wiki/Michael_Winslow
Michael Winterbottom	http://en.wikipedia.org/wiki/Michael_Winterbottom
Michael Yonkers	http://en.wikipedia.org/wiki/Michael_Yonkers
Michael York	http://en.wikipedia.org/wiki/Michael_York_(actor)
Micha�lle Jean	http://en.wikipedia.org/wiki/Micha%EBlle_Jean
Michel de Castelnau	http://en.wikipedia.org/wiki/Michel_de_Castelnau
Michel de Ghelderode	http://en.wikipedia.org/wiki/Michel_de_Ghelderode
Michel de Montaigne	http://en.wikipedia.org/wiki/Michel_de_Montaigne
Michel Foucault	http://en.wikipedia.org/wiki/Michel_Foucault
Michel Gondry	http://en.wikipedia.org/wiki/Michel_Gondry
Michel Legrand	http://en.wikipedia.org/wiki/Michel_Legrand
Michel Magne	http://en.wikipedia.org/wiki/Michel_Magne
Michel Mathieu	http://en.wikipedia.org/wiki/Michel_Mathieu
Michel Ney	http://en.wikipedia.org/wiki/Michel_Ney
Michel Platini	http://en.wikipedia.org/wiki/Michel_Platini
Michel Roger	http://en.wikipedia.org/wiki/Michel_Roger
Michel Suleiman	http://en.wikipedia.org/wiki/Michel_Suleiman
Michelangelo Antonioni	http://en.wikipedia.org/wiki/Michelangelo_Antonioni
Michele Bachmann	http://en.wikipedia.org/wiki/Michele_Bachmann
Michele Lee	http://en.wikipedia.org/wiki/Michele_Lee
Mich�le Mercier	http://en.wikipedia.org/wiki/Mich%E8le_Mercier
Mich�le Morgan	http://en.wikipedia.org/wiki/Mich%E8le_Morgan
Michel-Eug�ne Chevreul	http://en.wikipedia.org/wiki/Michel-Eug%E8ne_Chevreul
Michelle Bachelet	http://en.wikipedia.org/wiki/Michelle_Bachelet
Michelle Bachelet	http://en.wikipedia.org/wiki/Michelle_Bachelet
Michelle Bernard	http://en.wikipedia.org/wiki/Michelle_Bernard
Michelle Branch	http://en.wikipedia.org/wiki/Michelle_Branch
Michelle Clunie	http://en.wikipedia.org/wiki/Michelle_Clunie
Michelle Gildernew	http://en.wikipedia.org/wiki/Michelle_Gildernew
Michelle Johnson	http://en.wikipedia.org/wiki/Michelle_Johnson_(actress)
Michelle Kwan	http://en.wikipedia.org/wiki/Michelle_Kwan
Michelle Leslie	http://en.wikipedia.org/wiki/Michelle_Leslie
Michelle Malkin	http://en.wikipedia.org/wiki/Michelle_Malkin
Michelle Malone	http://en.wikipedia.org/wiki/Michelle_Malone
Michelle Pfeiffer	http://en.wikipedia.org/wiki/Michelle_Pfeiffer
Michelle Phillips	http://en.wikipedia.org/wiki/Michelle_Phillips
Michelle Rodriguez	http://en.wikipedia.org/wiki/Michelle_Rodriguez
Michelle Shocked	http://en.wikipedia.org/wiki/Michelle_Shocked
Michelle Thomas	http://en.wikipedia.org/wiki/Michelle_Thomas
Michelle Trachtenberg	http://en.wikipedia.org/wiki/Michelle_Trachtenberg
Michelle Wie	http://en.wikipedia.org/wiki/Michelle_Wie
Michelle Williams	http://en.wikipedia.org/wiki/Michelle_Williams_(actress)
Michelle Williams	http://en.wikipedia.org/wiki/Michelle_Williams_(singer)
Michelle Yeoh	http://en.wikipedia.org/wiki/Michelle_Yeoh
Michiko Kakutani	http://en.wikipedia.org/wiki/Michiko_Kakutani
Mick Avory	http://en.wikipedia.org/wiki/Mick_Avory
Mick Fleetwood	http://en.wikipedia.org/wiki/Mick_Fleetwood
Mick Foley	http://en.wikipedia.org/wiki/Mick_Foley
Mick Jagger	http://en.wikipedia.org/wiki/Mick_Jagger
Mick Jones	http://en.wikipedia.org/wiki/Mick_Jones_(singer,_born_1944)
Mick Jones	http://en.wikipedia.org/wiki/Mick_Jones_(The_Clash)
Mick Mars	http://en.wikipedia.org/wiki/Mick_Mars
Mick Ralphs	http://en.wikipedia.org/wiki/Mick_Ralphs
Mick Ronson	http://en.wikipedia.org/wiki/Mick_Ronson
Mick Taylor	http://en.wikipedia.org/wiki/Mick_Taylor
Mickey Cochrane	http://en.wikipedia.org/wiki/Mickey_Cochrane
Mickey Edwards	http://en.wikipedia.org/wiki/Mickey_Edwards
Mickey Gilley	http://en.wikipedia.org/wiki/Mickey_Gilley
Mickey Hart	http://en.wikipedia.org/wiki/Mickey_Hart
Mickey Kantor	http://en.wikipedia.org/wiki/Mickey_Kantor
Mickey Leland	http://en.wikipedia.org/wiki/Mickey_Leland
Mickey Mantle	http://en.wikipedia.org/wiki/Mickey_Mantle
Mickey Rooney	http://en.wikipedia.org/wiki/Mickey_Rooney
Mickey Rourke	http://en.wikipedia.org/wiki/Mickey_Rourke
Mickey Spillane	http://en.wikipedia.org/wiki/Mickey_Spillane
Micky Dolenz	http://en.wikipedia.org/wiki/Micky_Dolenz
Midge Decter	http://en.wikipedia.org/wiki/Midge_Decter
Midge Ure	http://en.wikipedia.org/wiki/Midge_Ure
Miguel Abia Biteo Borico	http://en.wikipedia.org/wiki/Miguel_Abia_Biteo_Borico
Miguel �ngel Asturias	http://en.wikipedia.org/wiki/Miguel_%C1ngel_Asturias
Miguel Bos�	http://en.wikipedia.org/wiki/Miguel_Bos%E9
Miguel Cabrera	http://en.wikipedia.org/wiki/Miguel_Cabrera
Miguel de Bragan�a	http://en.wikipedia.org/wiki/Miguel_de_Bragan%C3%A7a
Miguel de Cervantes	http://en.wikipedia.org/wiki/Miguel_de_Cervantes
Miguel de Icaza	http://en.wikipedia.org/wiki/Miguel_de_Icaza
Miguel de Unamuno	http://en.wikipedia.org/wiki/Miguel_de_Unamuno
Miguel Ferrer	http://en.wikipedia.org/wiki/Miguel_Ferrer
Miguel Hern�ndez	http://en.wikipedia.org/wiki/Miguel_Hern%E1ndez
Miguel Hidalgo	http://en.wikipedia.org/wiki/Miguel_Hidalgo
Miguel Sandoval	http://en.wikipedia.org/wiki/Miguel_Sandoval
Mihai Eminescu	http://en.wikipedia.org/wiki/Mihai_Eminescu
Mih�ly Csokonai Vit�z	http://en.wikipedia.org/wiki/Mih%E1ly_Csokonai_Vit%E9z
Miho Hatori	http://en.wikipedia.org/wiki/Miho_Hatori
Mijailo Mijailovic	http://en.wikipedia.org/wiki/Mijailo_Mijailovic
Mika Boorem	http://en.wikipedia.org/wiki/Mika_Boorem
Mika H�kkinen	http://en.wikipedia.org/wiki/Mika_H%E4kkinen
Mike Allen	http://en.wikipedia.org/wiki/Michael_Allen_(journalist)
Mike Allsup	http://en.wikipedia.org/wiki/Mike_Allsup
Mike Aulby	http://en.wikipedia.org/wiki/Mike_Aulby
Mike Bibby	http://en.wikipedia.org/wiki/Mike_Bibby
Mike Bloomfield	http://en.wikipedia.org/wiki/Mike_Bloomfield
Mike Castle	http://en.wikipedia.org/wiki/Mike_Castle
Mike Coffman	http://en.wikipedia.org/wiki/Mike_Coffman
Mike Conaway	http://en.wikipedia.org/wiki/Mike_Conaway
Mike Connors	http://en.wikipedia.org/wiki/Mike_Connors
Mike Crockart	http://en.wikipedia.org/wiki/Mike_Crockart
Mike Curb	http://en.wikipedia.org/wiki/Mike_Curb
Mike D	http://en.wikipedia.org/wiki/Mike_D
Mike DeWine	http://en.wikipedia.org/wiki/Mike_DeWine
Mike Diana	http://en.wikipedia.org/wiki/Mike_Diana
Mike Dirnt	http://en.wikipedia.org/wiki/Mike_Dirnt
Mike Ditka	http://en.wikipedia.org/wiki/Mike_Ditka
Mike Douglas	http://en.wikipedia.org/wiki/Mike_Douglas
Mike Doyle	http://en.wikipedia.org/wiki/Michael_F._Doyle
Mike Easley	http://en.wikipedia.org/wiki/Mike_Easley
Mike Epps	http://en.wikipedia.org/wiki/Mike_Epps
Mike Espy	http://en.wikipedia.org/wiki/Mike_Espy
Mike Farrell	http://en.wikipedia.org/wiki/Mike_Farrell
Mike Figgis	http://en.wikipedia.org/wiki/Mike_Figgis
Mike Fitzpatrick	http://en.wikipedia.org/wiki/Mike_Fitzpatrick
Mike Freer	http://en.wikipedia.org/wiki/Mike_Freer
Mike Gallagher	http://en.wikipedia.org/wiki/Mike_Gallagher
Mike Gapes	http://en.wikipedia.org/wiki/Mike_Gapes
Mike Gordon	http://en.wikipedia.org/wiki/Mike_Gordon
Mike Gravel	http://en.wikipedia.org/wiki/Mike_Gravel
Mike Hancock	http://en.wikipedia.org/wiki/Mike_Hancock_(UK_politician)
Mike Honda	http://en.wikipedia.org/wiki/Mike_Honda
Mike Huckabee	http://en.wikipedia.org/wiki/Mike_Huckabee
Mike Huckabee	http://en.wikipedia.org/wiki/Mike_Huckabee
Mike Johanns	http://en.wikipedia.org/wiki/Mike_Johanns
Mike Jones	http://en.wikipedia.org/wiki/Mike_Jones_(rapper)
Mike Judge	http://en.wikipedia.org/wiki/Mike_Judge
Mike Leigh	http://en.wikipedia.org/wiki/Mike_Leigh
Mike Lookinland	http://en.wikipedia.org/wiki/Mike_Lookinland
Mike Love	http://en.wikipedia.org/wiki/Mike_Love
Mike Lowry	http://en.wikipedia.org/wiki/Mike_Lowry
Mike Mansfield	http://en.wikipedia.org/wiki/Mike_Mansfield
Mike McCready	http://en.wikipedia.org/wiki/Mike_McCready
Mike McCurry	http://en.wikipedia.org/wiki/Mike_McCurry_(press_secretary)
Mike McIntyre	http://en.wikipedia.org/wiki/Mike_McIntyre
Mike Mills	http://en.wikipedia.org/wiki/Mike_Mills
Mike Myers	http://en.wikipedia.org/wiki/Mike_Myers_(actor)
Mike Nesmith	http://en.wikipedia.org/wiki/Mike_Nesmith
Mike Ness	http://en.wikipedia.org/wiki/Mike_Ness
Mike Newell	http://en.wikipedia.org/wiki/Mike_Newell_(director)
Mike Nichols	http://en.wikipedia.org/wiki/Mike_Nichols
Mike O'Callaghan	http://en.wikipedia.org/wiki/Mike_O%27Callaghan
Mike Oldfield	http://en.wikipedia.org/wiki/Mike_Oldfield
Mike O'Malley	http://en.wikipedia.org/wiki/Mike_O%27Malley
Mike Paradinas	http://en.wikipedia.org/wiki/Mike_Paradinas
Mike Patton	http://en.wikipedia.org/wiki/Mike_Patton
Mike Pence	http://en.wikipedia.org/wiki/Mike_Pence
Mike Penning	http://en.wikipedia.org/wiki/Mike_Penning
Mike Peters	http://en.wikipedia.org/wiki/Mike_Peters_(musician)
Mike Piazza	http://en.wikipedia.org/wiki/Mike_Piazza
Mike Portnoy	http://en.wikipedia.org/wiki/Mike_Portnoy
Mike Ratledge	http://en.wikipedia.org/wiki/Mike_Ratledge
Mike Rogers	http://en.wikipedia.org/wiki/Mike_D._Rogers
Mike Rogers	http://en.wikipedia.org/wiki/Mike_Rogers_(Michigan_politician)
Mike Ross	http://en.wikipedia.org/wiki/Mike_Ross
Mike Rounds	http://en.wikipedia.org/wiki/Mike_Rounds
Mike Royko	http://en.wikipedia.org/wiki/Mike_Royko
Mike Rozier	http://en.wikipedia.org/wiki/Mike_Rozier
Mike Rutherford	http://en.wikipedia.org/wiki/Mike_Rutherford
Mike Schmidt	http://en.wikipedia.org/wiki/Mike_Schmidt
Mike Shinoda	http://en.wikipedia.org/wiki/Mike_Shinoda
Mike Simpson	http://en.wikipedia.org/wiki/Mike_Simpson
Mike Singletary	http://en.wikipedia.org/wiki/Mike_Singletary
Mike Sodrel	http://en.wikipedia.org/wiki/Mike_Sodrel
Mike Stoller	http://en.wikipedia.org/wiki/Mike_Stoller
Mike Straka	http://en.wikipedia.org/wiki/Mike_Straka
Mike Strang	http://en.wikipedia.org/wiki/Mike_Strang
Mike Synar	http://en.wikipedia.org/wiki/Mike_Synar
Mike Thompson	http://en.wikipedia.org/wiki/Mike_Thompson
Mike Tyson	http://en.wikipedia.org/wiki/Mike_Tyson
Mike Vogel	http://en.wikipedia.org/wiki/Mike_Vogel
Mike Wallace	http://en.wikipedia.org/wiki/Mike_Wallace_(journalist)
Mike Watt	http://en.wikipedia.org/wiki/Mike_Watt
Mike Weatherley	http://en.wikipedia.org/wiki/Mike_Weatherley
Mike Weir	http://en.wikipedia.org/wiki/Mike_Weir_(SNP)
Mike Wilson	http://en.wikipedia.org/wiki/Mike_Wilson_(filmmaker)
Mike Wood	http://en.wikipedia.org/wiki/Mike_Wood_(politician)
Mikey Way	http://en.wikipedia.org/wiki/Mikey_Way
Mikhail An	http://en.wikipedia.org/wiki/Mikhail_An
Mikhail Bakunin	http://en.wikipedia.org/wiki/Mikhail_Bakunin
Mikhail Baryshnikov	http://en.wikipedia.org/wiki/Mikhail_Baryshnikov
Mikhail Bulgakov	http://en.wikipedia.org/wiki/Mikhail_Bulgakov
Mikhail Fradkov	http://en.wikipedia.org/wiki/Mikhail_Fradkov
Mikhail Fradkov	http://en.wikipedia.org/wiki/Mikhail_Fradkov
Mikhail Glinka	http://en.wikipedia.org/wiki/Mikhail_Glinka
Mikhail Gorbachev	http://en.wikipedia.org/wiki/Mikhail_Gorbachev
Mikhail Kasyanov	http://en.wikipedia.org/wiki/Mikhail_Kasyanov
Mikhail Khodorkovsky	http://en.wikipedia.org/wiki/Mikhail_Khodorkovsky
Mikhail Lermontov	http://en.wikipedia.org/wiki/Mikhail_Lermontov
Mikhail Lomonosov	http://en.wikipedia.org/wiki/Mikhail_Lomonosov
Mikhail Saakashvili	http://en.wikipedia.org/wiki/Mikhail_Saakashvili
Mikhail Saakashvili	http://en.wikipedia.org/wiki/Mikhail_Saakashvili
Mikhail Timofeyevich Kalashnikov	http://en.wikipedia.org/wiki/Mikhail_Kalashnikov
Mikheil Saakashvili	http://en.wikipedia.org/wiki/Mikheil_Saakashvili
Miki Berenyi	http://en.wikipedia.org/wiki/Miki_Berenyi
Mikul� Dzurinda	http://en.wikipedia.org/wiki/Mikul%E1%9A_Dzurinda
Mila Kunis	http://en.wikipedia.org/wiki/Mila_Kunis
Milan Kundera	http://en.wikipedia.org/wiki/Milan_Kundera
Milburn Stone	http://en.wikipedia.org/wiki/Milburn_Stone
Mildred Wirt Benson	http://en.wikipedia.org/wiki/Mildred_Wirt_Benson
Miles Ambrose	http://en.wikipedia.org/wiki/Miles_Ambrose
Miles Copeland	http://en.wikipedia.org/wiki/Miles_Copeland
Miles D. White	http://en.wikipedia.org/wiki/Miles_D._White
Miles Davis	http://en.wikipedia.org/wiki/Miles_Davis
Miles Poindexter	http://en.wikipedia.org/wiki/Miles_Poindexter
Milla Jovovich	http://en.wikipedia.org/wiki/Milla_Jovovich
Millard E. Tydings	http://en.wikipedia.org/wiki/Millard_E._Tydings
Millard Fillmore	http://en.wikipedia.org/wiki/Millard_Fillmore
Milo �ukanovic	http://en.wikipedia.org/wiki/Milo_Đukanović
Milo Ventimiglia	http://en.wikipedia.org/wiki/Milo_Ventimiglia
Milorad Dodik	http://en.wikipedia.org/wiki/Milorad_Dodik
Milos Forman	http://en.wikipedia.org/wiki/Milos_Forman
Milton Babbitt	http://en.wikipedia.org/wiki/Milton_Babbitt
Milton Berle	http://en.wikipedia.org/wiki/Milton_Berle
Milton Friedman	http://en.wikipedia.org/wiki/Milton_Friedman
Milton Obote	http://en.wikipedia.org/wiki/Milton_Obote
Milton Sills	http://en.wikipedia.org/wiki/Milton_Sills
Mily Balakirev	http://en.wikipedia.org/wiki/Mily_Balakirev
Mimi Rogers	http://en.wikipedia.org/wiki/Mimi_Rogers
Mindy Cohn	http://en.wikipedia.org/wiki/Mindy_Cohn
Mindy McCready	http://en.wikipedia.org/wiki/Mindy_McCready
Ming Yao	http://en.wikipedia.org/wiki/Ming_Yao
Mink Stole	http://en.wikipedia.org/wiki/Mink_Stole
Minna Aaltonen	http://en.wikipedia.org/wiki/Minna_Aaltonen
Minnesota Fats	http://en.wikipedia.org/wiki/Rudolf_Wanderone
Minnie Driver	http://en.wikipedia.org/wiki/Minnie_Driver
Minnie Pearl	http://en.wikipedia.org/wiki/Minnie_Pearl
Mir Aimal Kasi	http://en.wikipedia.org/wiki/Mir_Aimal_Kasi
Mira Calix	http://en.wikipedia.org/wiki/Mira_Calix
Mira Nair	http://en.wikipedia.org/wiki/Mira_Nair
Mira Sorvino	http://en.wikipedia.org/wiki/Mira_Sorvino
Miranda Otto	http://en.wikipedia.org/wiki/Miranda_Otto
Miranda Richardson	http://en.wikipedia.org/wiki/Miranda_Richardson
Mircea Albulescu	http://en.wikipedia.org/wiki/Mircea_Albulescu
Mireille Mathieu	http://en.wikipedia.org/wiki/Mireille_Mathieu
Miriam Hopkins	http://en.wikipedia.org/wiki/Miriam_Hopkins
Mirko Cvetkovic	http://en.wikipedia.org/wiki/Mirko_Cvetkovic
Mischa Auer	http://en.wikipedia.org/wiki/Mischa_Auer
Mischa Barton	http://en.wikipedia.org/wiki/Mischa_Barton
Miss Cleo	http://en.wikipedia.org/wiki/Miss_Cleo
Missy Elliott	http://en.wikipedia.org/wiki/Missy_Elliott
Missy Gold	http://en.wikipedia.org/wiki/Missy_Gold
Missy Higgins	http://en.wikipedia.org/wiki/Missy_Higgins
Misty Mundae	http://en.wikipedia.org/wiki/Misty_Mundae
Mitch Albom	http://en.wikipedia.org/wiki/Mitch_Albom
Mitch Daniels	http://en.wikipedia.org/wiki/Mitch_Daniels
Mitch Daniels	http://en.wikipedia.org/wiki/Mitch_Daniels
Mitch Hedberg	http://en.wikipedia.org/wiki/Mitch_Hedberg
Mitch Kapor	http://en.wikipedia.org/wiki/Mitch_Kapor
Mitch Landrieu	http://en.wikipedia.org/wiki/Mitch_Landrieu
Mitch McConnell	http://en.wikipedia.org/wiki/Mitch_McConnell
Mitch McConnell	http://en.wikipedia.org/wiki/Mitch_McConnell
Mitch Miller	http://en.wikipedia.org/wiki/Mitch_Miller
Mitch Mitchell	http://en.wikipedia.org/wiki/Mitch_Mitchell
Mitch Pileggi	http://en.wikipedia.org/wiki/Mitch_Pileggi
Mitt Romney	http://en.wikipedia.org/wiki/Mitt_Romney
Mitzi Gaynor	http://en.wikipedia.org/wiki/Mitzi_Gaynor
Mitzi Kapture	http://en.wikipedia.org/wiki/Mitzi_Kapture
Miyamoto Musashi	http://en.wikipedia.org/wiki/Miyamoto_Musashi
Miyeegombo Enkhbold	http://en.wikipedia.org/wiki/Miyeegombo_Enkhbold
Miyoshi Umeki	http://en.wikipedia.org/wiki/Miyoshi_Umeki
Mizan Zainal Abidin	http://en.wikipedia.org/wiki/Mizan_Zainal_Abidin
Mizengo Pinda	http://en.wikipedia.org/wiki/Mizengo_Pinda
Mo Collins	http://en.wikipedia.org/wiki/Mo_Collins
Mo Rocca	http://en.wikipedia.org/wiki/Mo_Rocca
Mo Udall	http://en.wikipedia.org/wiki/Mo_Udall
Mobutu Sese Seko	http://en.wikipedia.org/wiki/Mobutu_Sese_Seko
Moby	http://en.wikipedia.org/wiki/Moby
Modest Mussorgsky	http://en.wikipedia.org/wiki/Modest_Mussorgsky
Modibo Sidib�	http://en.wikipedia.org/wiki/Modibo_Sidib%E9
Moe Howard	http://en.wikipedia.org/wiki/Moe_Howard
Mohamed Abdul Quasim al-Zwai	http://en.wikipedia.org/wiki/Mohamed_Abdul_Quasim_al-Zwai
Mohamed al-Fayed	http://en.wikipedia.org/wiki/Mohamed_al-Fayed
Mohamed al-Otari	http://en.wikipedia.org/wiki/Muhammad_Naji_al-Otari
Mohamed Bacar	http://en.wikipedia.org/wiki/Mohamed_Bacar
Mohamed El Baradei	http://en.wikipedia.org/wiki/Mohamed_El_Baradei
Mohamed Ghannouchi	http://en.wikipedia.org/wiki/Mohamed_Ghannouchi
Mohamed Nasheed	http://en.wikipedia.org/wiki/Mohamed_Nasheed
Mohamed Ould Abdel Aziz	http://en.wikipedia.org/wiki/Mohamed_Ould_Abdel_Aziz
Mohamed Said Fazul	http://en.wikipedia.org/wiki/Mohamed_Said_Fazul
Mohammad Ali Jinnah	http://en.wikipedia.org/wiki/Mohammad_Ali_Jinnah
Mohammad Khatami	http://en.wikipedia.org/wiki/Mohammad_Khatami
Mohammad Najibullah	http://en.wikipedia.org/wiki/Mohammad_Najibullah
Mohammad Rabbani	http://en.wikipedia.org/wiki/Mohammad_Rabbani
Mohammed Abdel Aziz	http://en.wikipedia.org/wiki/Mohammed_Abdel_Aziz
Mohammed Atta	http://en.wikipedia.org/wiki/Mohammed_Atta
Mohammed bin Rashid Al Maktoum	http://en.wikipedia.org/wiki/Mohammed_bin_Rashid_Al_Maktoum
Mohammed Jamal Khalifa	http://en.wikipedia.org/wiki/Mohammed_Jamal_Khalifa
Mohammed Omar	http://en.wikipedia.org/wiki/Mohammed_Omar
Mohammed VI	http://en.wikipedia.org/wiki/Mohammed_VI
Mohamud Muse Hersi "Adde"	http://en.wikipedia.org/wiki/Mohamud_Muse_Hersi
Mohandas Ghandi	http://en.wikipedia.org/wiki/Mohandas_Ghandi
Moira Kelly	http://en.wikipedia.org/wiki/Moira_Kelly
Moira Shearer	http://en.wikipedia.org/wiki/Moira_Shearer
Moise Tshombe	http://en.wikipedia.org/wiki/Moise_Tshombe
Mojo Nixon	http://en.wikipedia.org/wiki/Mojo_Nixon
Mollie Sugden	http://en.wikipedia.org/wiki/Mollie_Sugden
Molly Ivins	http://en.wikipedia.org/wiki/Molly_Ivins
Molly Parker	http://en.wikipedia.org/wiki/Molly_Parker
Molly Price	http://en.wikipedia.org/wiki/Molly_Price
Molly Ringwald	http://en.wikipedia.org/wiki/Molly_Ringwald
Molly Shannon	http://en.wikipedia.org/wiki/Molly_Shannon
Molly Sims	http://en.wikipedia.org/wiki/Molly_Sims
Molly Yard	http://en.wikipedia.org/wiki/Molly_Yard
Mona Charen	http://en.wikipedia.org/wiki/Mona_Charen
Mona Van Duyn	http://en.wikipedia.org/wiki/Mona_Van_Duyn
Mongo Santamaria	http://en.wikipedia.org/wiki/Mongo_Santamaria
Monica Bellucci	http://en.wikipedia.org/wiki/Monica_Bellucci
Monica Crowley	http://en.wikipedia.org/wiki/Monica_Crowley
Monica Keena	http://en.wikipedia.org/wiki/Monica_Keena
Monica Lewinsky	http://en.wikipedia.org/wiki/Monica_Lewinsky
Monica Potter	http://en.wikipedia.org/wiki/Monica_Potter
Monica Seles	http://en.wikipedia.org/wiki/Monica_Seles
Moniza Alvi	http://en.wikipedia.org/wiki/Moniza_Alvi
Monte Blue	http://en.wikipedia.org/wiki/Monte_Blue
Montel Williams	http://en.wikipedia.org/wiki/Montel_Williams
Montezuma II	http://en.wikipedia.org/wiki/Montezuma_II
Montgomery Clift	http://en.wikipedia.org/wiki/Montgomery_Clift
Monty Hall	http://en.wikipedia.org/wiki/Monty_Hall
Monty Woolley	http://en.wikipedia.org/wiki/Monty_Woolley
Moon Unit Zappa	http://en.wikipedia.org/wiki/Moon_Unit_Zappa
Morarji Desai	http://en.wikipedia.org/wiki/Morarji_Desai
Mordecai Brown	http://en.wikipedia.org/wiki/Mordecai_Brown
Mordecai Richler	http://en.wikipedia.org/wiki/Mordecai_Richler
Mordechai Vanunu	http://en.wikipedia.org/wiki/Mordechai_Vanunu
Morey Amsterdam	http://en.wikipedia.org/wiki/Morey_Amsterdam
Morgan Alling	http://en.wikipedia.org/wiki/Morgan_Alling
Morgan Brittany	http://en.wikipedia.org/wiki/Morgan_Brittany
Morgan Fairchild	http://en.wikipedia.org/wiki/Morgan_Fairchild
Morgan Freeman	http://en.wikipedia.org/wiki/Morgan_Freeman
Morgan Lewis	http://en.wikipedia.org/wiki/Morgan_Lewis_(governor)
Morgan Spurlock	http://en.wikipedia.org/wiki/Morgan_Spurlock
Morgan Tsvangirai	http://en.wikipedia.org/wiki/Morgan_Tsvangirai
Morgan Woodward	http://en.wikipedia.org/wiki/Morgan_Woodward
Moritz Hartmann	http://en.wikipedia.org/wiki/Moritz_Hartmann
Moritz Leuenberger	http://en.wikipedia.org/wiki/Moritz_Leuenberger
Moritz Schlick	http://en.wikipedia.org/wiki/Moritz_Schlick
Morley Callaghan	http://en.wikipedia.org/wiki/Morley_Callaghan
Morley Safer	http://en.wikipedia.org/wiki/Morley_Safer
Morris Chestnut	http://en.wikipedia.org/wiki/Morris_Chestnut
Morris Day	http://en.wikipedia.org/wiki/Morris_Day
Morris Dees	http://en.wikipedia.org/wiki/Morris_Dees
Morris K. Udall	http://en.wikipedia.org/wiki/Morris_K._Udall
Morris Louis	http://en.wikipedia.org/wiki/Morris_Louis
Morrison Waite	http://en.wikipedia.org/wiki/Morrison_Waite
Morrissey	http://en.wikipedia.org/wiki/Morrissey
Mort Kondracke	http://en.wikipedia.org/wiki/Mort_Kondracke
Mort Sahl	http://en.wikipedia.org/wiki/Mort_Sahl
Mort Zuckerman	http://en.wikipedia.org/wiki/Mort_Zuckerman
Mortimer J. Adler	http://en.wikipedia.org/wiki/Mortimer_J._Adler
Mortimer Wheeler	http://en.wikipedia.org/wiki/Mortimer_Wheeler
Morton C. Blackwell	http://en.wikipedia.org/wiki/Morton_C._Blackwell
Morton Downey, Jr.	http://en.wikipedia.org/wiki/Morton_Downey%2C_Jr.
Morton Feldman	http://en.wikipedia.org/wiki/Morton_Feldman
Morton Heilig	http://en.wikipedia.org/wiki/Morton_Heilig
Morton Stevens	http://en.wikipedia.org/wiki/Morton_Stevens
Mos Def	http://en.wikipedia.org/wiki/Mos_Def
Mose Allison	http://en.wikipedia.org/wiki/Mose_Allison
Moses de Leon	http://en.wikipedia.org/wiki/Moses_de_Leon
Moses Malone	http://en.wikipedia.org/wiki/Moses_Malone
Moses Mendelssohn	http://en.wikipedia.org/wiki/Moses_Mendelssohn
Moses Sithole	http://en.wikipedia.org/wiki/Moses_Sithole
Moshe Dayan	http://en.wikipedia.org/wiki/Moshe_Dayan
Moshe Katsav	http://en.wikipedia.org/wiki/Moshe_Katsav
Moshe Katsav	http://en.wikipedia.org/wiki/Moshe_Katsav
Moshe Sharett	http://en.wikipedia.org/wiki/Moshe_Sharett
Moss Hart	http://en.wikipedia.org/wiki/Moss_Hart
Mossimo Giannulli	http://en.wikipedia.org/wiki/Mossimo_Giannulli
Mother Angelica	http://en.wikipedia.org/wiki/Mother_Angelica
Mother Shipton	http://en.wikipedia.org/wiki/Mother_Shipton
Mother Teresa	http://en.wikipedia.org/wiki/Mother_Teresa
Moulaye Ould Mohamed Laghdaf	http://en.wikipedia.org/wiki/Moulaye_Ould_Mohamed_Laghdaf
Mounir el-Motassadeq	http://en.wikipedia.org/wiki/Mounir_el-Motassadeq
Moussa Dadis Camara	http://en.wikipedia.org/wiki/Moussa_Dadis_Camara
Moustapha Akkad	http://en.wikipedia.org/wiki/Moustapha_Akkad
Mr. Blackwell	http://en.wikipedia.org/wiki/Mr._Blackwell
Mr. Lif	http://en.wikipedia.org/wiki/Mr._Lif
Mr. T	http://en.wikipedia.org/wiki/Mr._T
Ms. Dynamite	http://en.wikipedia.org/wiki/Ms._Dynamite
Ms. Jade	http://en.wikipedia.org/wiki/Ms._Jade
Mswati III	http://en.wikipedia.org/wiki/Mswati_III
Muammar al-Gaddafi	http://en.wikipedia.org/wiki/Muammar_al-Gaddafi
Muddy Waters	http://en.wikipedia.org/wiki/Muddy_Waters
Muhal Richard Abrams	http://en.wikipedia.org/wiki/Muhal_Richard_Abrams
Muhammad Ali	http://en.wikipedia.org/wiki/Muhammad_Ali
Muhammad al-Otari	http://en.wikipedia.org/wiki/Muhammad_al-Otari
Muhammad Yunus	http://en.wikipedia.org/wiki/Muhammad_Yunus
Muhammad Zia-ul-Haq	http://en.wikipedia.org/wiki/Muhammad_Zia-ul-Haq
Muhammed Saeed al-Sahaf	http://en.wikipedia.org/wiki/Muhammed_Saeed_al-Sahaf
Mujibur Rahman	http://en.wikipedia.org/wiki/Mujibur_Rahman
Mukesh Ambani	http://en.wikipedia.org/wiki/Mukesh_Ambani
Mulk Raj Anand	http://en.wikipedia.org/wiki/Mulk_Raj_Anand
Mumia Abu-Jamal	http://en.wikipedia.org/wiki/Mumia_Abu-Jamal
Mungo Park	http://en.wikipedia.org/wiki/Mungo_Park_(explorer)
Munro Leaf	http://en.wikipedia.org/wiki/Munro_Leaf
Muqtada al-Sadr	http://en.wikipedia.org/wiki/Muqtada_al-Sadr
Murad I	http://en.wikipedia.org/wiki/Murad_I
Murad II	http://en.wikipedia.org/wiki/Murad_II
Muriel Aked	http://en.wikipedia.org/wiki/Muriel_Aked
Muriel Rukeyser	http://en.wikipedia.org/wiki/Muriel_Rukeyser
Muriel Spark	http://en.wikipedia.org/wiki/Muriel_Spark
Murray Gell-Mann	http://en.wikipedia.org/wiki/Murray_Gell-Mann
Murray Head	http://en.wikipedia.org/wiki/Murray_Head
Murray Krieger	http://en.wikipedia.org/wiki/Murray_Krieger
Murray Rose	http://en.wikipedia.org/wiki/Murray_Rose
Murray Rothbard	http://en.wikipedia.org/wiki/Murray_Rothbard
Murray Waas	http://en.wikipedia.org/wiki/Murray_Waas
Mushroom	http://en.wikipedia.org/wiki/Andrew_Vowles
Mustafa Altioklar	http://en.wikipedia.org/wiki/Mustafa_Altioklar
Mustapha Adouani	http://en.wikipedia.org/wiki/Mustapha_Adouani
Mutt Lange	http://en.wikipedia.org/wiki/Mutt_Lange
Muttiah Muralitharan	http://en.wikipedia.org/wiki/Muttiah_Muralitharan
Muzio Clementi	http://en.wikipedia.org/wiki/Muzio_Clementi
Mwai Kibaki	http://en.wikipedia.org/wiki/Mwai_Kibaki
Mya	http://en.wikipedia.org/wiki/Mýa
Mykola Azarov	http://en.wikipedia.org/wiki/Mykola_Azarov
Myra Hindley	http://en.wikipedia.org/wiki/Myra_Hindley
Myrna Blyth	http://en.wikipedia.org/wiki/Myrna_Blyth
Myrna Loy	http://en.wikipedia.org/wiki/Myrna_Loy
Myron C. Taylor	http://en.wikipedia.org/wiki/Myron_C._Taylor
Myron Floren	http://en.wikipedia.org/wiki/Myron_Floren
N. Scott Momaday	http://en.wikipedia.org/wiki/N._Scott_Momaday
Nabih Berri	http://en.wikipedia.org/wiki/Nabih_Berri
Nadhim Zahawi	http://en.wikipedia.org/wiki/Nadhim_Zahawi
Nadia Bjorlin	http://en.wikipedia.org/wiki/Nadia_Bjorlin
Nadia Comaneci	http://en.wikipedia.org/wiki/Nadia_Comaneci
Nadia Petrova	http://en.wikipedia.org/wiki/Nadia_Petrova
Nadine Dorries	http://en.wikipedia.org/wiki/Nadine_Dorries
Nadine Gordimer	http://en.wikipedia.org/wiki/Nadine_Gordimer
Nafisa Joseph	http://en.wikipedia.org/wiki/Nafisa_Joseph
Naguib Mahfouz	http://en.wikipedia.org/wiki/Naguib_Mahfouz
Nahas Angula	http://en.wikipedia.org/wiki/Nahas_Angula
Nahum Tate	http://en.wikipedia.org/wiki/Nahum_Tate
Naima Akef	http://en.wikipedia.org/wiki/Naima_Akef
Najib Razak	http://en.wikipedia.org/wiki/Najib_Razak
Nam June Paik	http://en.wikipedia.org/wiki/Nam_June_Paik
Nambaryn Enkhbayar	http://en.wikipedia.org/wiki/Nambaryn_Enkhbayar
Nan Kempner	http://en.wikipedia.org/wiki/Nan_Kempner
Nana Vasconcelos	http://en.wikipedia.org/wiki/Nana_Vasconcelos
Nana Visitor	http://en.wikipedia.org/wiki/Nana_Visitor
Nancy Addison	http://en.wikipedia.org/wiki/Nancy_Addison
Nancy Allen	http://en.wikipedia.org/wiki/Nancy_Allen_(actress)
Nancy Alvarez	http://en.wikipedia.org/wiki/Nancy_Alvarez_%28triathlete%29
Nancy Astor	http://en.wikipedia.org/wiki/Nancy_Astor
Nancy Cartwright	http://en.wikipedia.org/wiki/Nancy_Cartwright
Nancy Grace	http://en.wikipedia.org/wiki/Nancy_Grace
Nancy Johnson	http://en.wikipedia.org/wiki/Nancy_Johnson
Nancy Kassebaum	http://en.wikipedia.org/wiki/Nancy_Kassebaum
Nancy Kerrigan	http://en.wikipedia.org/wiki/Nancy_Kerrigan
Nancy Kulp	http://en.wikipedia.org/wiki/Nancy_Kulp
Nancy Kwan	http://en.wikipedia.org/wiki/Nancy_Kwan
Nancy L. Johnson	http://en.wikipedia.org/wiki/Nancy_L._Johnson
Nancy Landon Kassebaum	http://en.wikipedia.org/wiki/Nancy_Landon_Kassebaum
Nancy Lopez	http://en.wikipedia.org/wiki/Nancy_Lopez
Nancy Marchand	http://en.wikipedia.org/wiki/Nancy_Marchand
Nancy McKeon	http://en.wikipedia.org/wiki/Nancy_McKeon
Nancy Mitford	http://en.wikipedia.org/wiki/Nancy_Mitford
Nancy O'Dell	http://en.wikipedia.org/wiki/Nancy_O%27Dell
Nancy Olson	http://en.wikipedia.org/wiki/Nancy_Olson
Nancy Pelosi	http://en.wikipedia.org/wiki/Nancy_Pelosi
Nancy Reagan	http://en.wikipedia.org/wiki/Nancy_Reagan
Nancy Sinatra	http://en.wikipedia.org/wiki/Nancy_Sinatra
Nancy Spungen	http://en.wikipedia.org/wiki/Nancy_Spungen
Nancy Travis	http://en.wikipedia.org/wiki/Nancy_Travis
Nancy Walker	http://en.wikipedia.org/wiki/Nancy_Walker
Nancy Walls	http://en.wikipedia.org/wiki/Nancy_Walls
Nancy Wilson	http://en.wikipedia.org/wiki/Nancy_Wilson_(rock_musician)
Nancy Wilson	http://en.wikipedia.org/wiki/Nancy_Wilson_(jazz_singer)
Nanette Fabray	http://en.wikipedia.org/wiki/Nanette_Fabray
Nanette Newman	http://en.wikipedia.org/wiki/Nanette_Newman
Naomi Campbell	http://en.wikipedia.org/wiki/Naomi_Campbell
Naomi Judd	http://en.wikipedia.org/wiki/Naomi_Judd
Naomi Klein	http://en.wikipedia.org/wiki/Naomi_Klein
Naomi Long	http://en.wikipedia.org/wiki/Naomi_Long
Naomi Watts	http://en.wikipedia.org/wiki/Naomi_Watts
Naomi Wolf	http://en.wikipedia.org/wiki/Naomi_Wolf
Naoto Kan	http://en.wikipedia.org/wiki/Naoto_Kan
Napoleon Bonaparte	http://en.wikipedia.org/wiki/Napoleon_Bonaparte
Napoleon II	http://en.wikipedia.org/wiki/Napoleon_II
Napoleon III	http://en.wikipedia.org/wiki/Napoleon_III
Napper Tandy	http://en.wikipedia.org/wiki/Napper_Tandy
Narasimha Rao	http://en.wikipedia.org/wiki/P._V._Narasimha_Rao
Nasser Muhammad Al Ahmad Al Sabah	http://en.wikipedia.org/wiki/Nasser_Muhammad_Al_Ahmad_Al_Sabah
Nastassja Kinski	http://en.wikipedia.org/wiki/Nastassja_Kinski
Nastassja Kinski	http://en.wikipedia.org/wiki/Nastassja_Kinski
Nat Hentoff	http://en.wikipedia.org/wiki/Nat_Hentoff
Nat King Cole	http://en.wikipedia.org/wiki/Nat_King_Cole
Nat Turner	http://en.wikipedia.org/wiki/Nat_Turner
Natalia Ginzburg	http://en.wikipedia.org/wiki/Natalia_Ginzburg
Natalie Appleton	http://en.wikipedia.org/wiki/Natalie_Appleton
Natalie Cole	http://en.wikipedia.org/wiki/Natalie_Cole
Natalie Imbruglia	http://en.wikipedia.org/wiki/Natalie_Imbruglia
Natalie Maines	http://en.wikipedia.org/wiki/Natalie_Maines
Natalie Merchant	http://en.wikipedia.org/wiki/Natalie_Merchant
Natalie Portman	http://en.wikipedia.org/wiki/Natalie_Portman
Natalie Schafer	http://en.wikipedia.org/wiki/Natalie_Schafer
Natalie Wood	http://en.wikipedia.org/wiki/Natalie_Wood
Natan Altman	http://en.wikipedia.org/wiki/Natan_Altman
Natas Kaupas	http://en.wikipedia.org/wiki/Natas_Kaupas
Natascha Engel	http://en.wikipedia.org/wiki/Natascha_Engel
Natascha McElhone	http://en.wikipedia.org/wiki/Natascha_McElhone
Natasha Bedingfield	http://en.wikipedia.org/wiki/Natasha_Bedingfield
Natasha Henstridge	http://en.wikipedia.org/wiki/Natasha_Henstridge
Natasha Lyonne	http://en.wikipedia.org/wiki/Natasha_Lyonne
Natasha Richardson	http://en.wikipedia.org/wiki/Natasha_Richardson
Nate Berkus	http://en.wikipedia.org/wiki/Nate_Berkus
Nate Dogg	http://en.wikipedia.org/wiki/Nate_Dogg
Nathalie Sarraute	http://en.wikipedia.org/wiki/Nathalie_Sarraute
Nathan Bailey	http://en.wikipedia.org/wiki/Nathan_Bailey
Nathan Bedford Forrest	http://en.wikipedia.org/wiki/Nathan_Bedford_Forrest
Nathan Deal	http://en.wikipedia.org/wiki/Nathan_Deal
Nathan Fillion	http://en.wikipedia.org/wiki/Nathan_Fillion
Nathan Glazer	http://en.wikipedia.org/wiki/Nathan_Glazer
Nathan Hale	http://en.wikipedia.org/wiki/Nathan_Hale
Nathan Lane	http://en.wikipedia.org/wiki/Nathan_Lane
Nathan M. Pusey	http://en.wikipedia.org/wiki/Nathan_M._Pusey
Nathan S�derblom	http://en.wikipedia.org/wiki/Nathan_S%F6derblom
Nathanael Greene	http://en.wikipedia.org/wiki/Nathanael_Greene
Nathanael West	http://en.wikipedia.org/wiki/Nathanael_West
Nathaniel Bacon	http://en.wikipedia.org/wiki/Nathaniel_Bacon_(politician)
Nathaniel Bar-Jonah	http://en.wikipedia.org/wiki/Nathaniel_Bar-Jonah
Nathaniel Hawthorne	http://en.wikipedia.org/wiki/Nathaniel_Hawthorne
Nathaniel P. Banks	http://en.wikipedia.org/wiki/Nathaniel_P._Banks
Nathaniel Parker Willis	http://en.wikipedia.org/wiki/Nathaniel_Parker_Willis
Nathaniel Pitcher	http://en.wikipedia.org/wiki/Nathaniel_Pitcher
Nathaniel Waena	http://en.wikipedia.org/wiki/Nathaniel_Waena
Nathaniel Ward	http://en.wikipedia.org/wiki/Nathaniel_Ward
Nathuram Vinayak Godse	http://en.wikipedia.org/wiki/Nathuram_Vinayak_Godse
Naum Gabo	http://en.wikipedia.org/wiki/Naum_Gabo
Naunton Wayne	http://en.wikipedia.org/wiki/Naunton_Wayne
Naveen Andrews	http://en.wikipedia.org/wiki/Naveen_Andrews
Navin  Ramgoolam	http://en.wikipedia.org/wiki/Navin__Ramgoolam
Neal Cassady	http://en.wikipedia.org/wiki/Neal_Cassady
Neal Conan	http://en.wikipedia.org/wiki/Neal_Conan
Neal Gabler	http://en.wikipedia.org/wiki/Neal_Gabler
Neal McDonough	http://en.wikipedia.org/wiki/Neal_McDonough
Neal Schon	http://en.wikipedia.org/wiki/Neal_Schon
Neal Smith	http://en.wikipedia.org/wiki/Neal_Edward_Smith
Neal Stephenson	http://en.wikipedia.org/wiki/Neal_Stephenson
Ned Beatty	http://en.wikipedia.org/wiki/Ned_Beatty
Nehemiah Grew	http://en.wikipedia.org/wiki/Nehemiah_Grew
Neil Abercrombie	http://en.wikipedia.org/wiki/Neil_Abercrombie
Neil Armstrong	http://en.wikipedia.org/wiki/Neil_Armstrong
Neil Bush	http://en.wikipedia.org/wiki/Neil_Bush
Neil Carmichael	http://en.wikipedia.org/wiki/Neil_Carmichael_(Conservative_politician)
Neil Cavuto	http://en.wikipedia.org/wiki/Neil_Cavuto
Neil Diamond	http://en.wikipedia.org/wiki/Neil_Diamond
Neil Finn	http://en.wikipedia.org/wiki/Neil_Finn
Neil Gaiman	http://en.wikipedia.org/wiki/Neil_Gaiman
Neil Goldschmidt	http://en.wikipedia.org/wiki/Neil_Goldschmidt
Neil H. McElroy	http://en.wikipedia.org/wiki/Neil_H._McElroy
Neil Innes	http://en.wikipedia.org/wiki/Neil_Innes
Neil Jordan	http://en.wikipedia.org/wiki/Neil_Jordan
Neil LaBute	http://en.wikipedia.org/wiki/Neil_LaBute
Neil Parish	http://en.wikipedia.org/wiki/Neil_Parish
Neil Patrick Harris	http://en.wikipedia.org/wiki/Neil_Patrick_Harris
Neil Peart	http://en.wikipedia.org/wiki/Neil_Peart
Neil Rudenstine	http://en.wikipedia.org/wiki/Neil_Rudenstine
Neil Sedaka	http://en.wikipedia.org/wiki/Neil_Sedaka
Neil Sheehan	http://en.wikipedia.org/wiki/Neil_Sheehan
Neil Simon	http://en.wikipedia.org/wiki/Neil_Simon
Neil Tennant	http://en.wikipedia.org/wiki/Neil_Tennant
Neil Walter	http://en.wikipedia.org/wiki/Neil_Walter
Neil Young	http://en.wikipedia.org/wiki/Neil_Young
Neko Case	http://en.wikipedia.org/wiki/Neko_Case
Nell Carter	http://en.wikipedia.org/wiki/Nell_Carter
Nella Larsen	http://en.wikipedia.org/wiki/Nella_Larsen
Nellie McKay	http://en.wikipedia.org/wiki/Nellie_McKay
Nelly Furtado	http://en.wikipedia.org/wiki/Nelly_Furtado
Nelson Algren	http://en.wikipedia.org/wiki/Nelson_Algren
Nelson Ascencio	http://en.wikipedia.org/wiki/Nelson_Ascencio
Nelson Bunker Hunt	http://en.wikipedia.org/wiki/Nelson_Bunker_Hunt
Nelson Burton, Jr.	http://en.wikipedia.org/wiki/Nelson_Burton%2C_Jr.
Nelson Dingley, Jr.	http://en.wikipedia.org/wiki/Nelson_Dingley%2C_Jr.
Nelson Eddy	http://en.wikipedia.org/wiki/Nelson_Eddy
Nelson Goodman	http://en.wikipedia.org/wiki/Nelson_Goodman
Nelson Mandela	http://en.wikipedia.org/wiki/Nelson_Mandela
Nelson O. Oduber	http://en.wikipedia.org/wiki/Nelson_O._Oduber
Nelson Rockefeller	http://en.wikipedia.org/wiki/Nelson_Rockefeller
Nelson W. Aldrich	http://en.wikipedia.org/wiki/Nelson_W._Aldrich
Neneh Cherry	http://en.wikipedia.org/wiki/Neneh_Cherry
N�stor Kirchner	http://en.wikipedia.org/wiki/N%E9stor_Kirchner
N�stor Kirchner	http://en.wikipedia.org/wiki/N%E9stor_Kirchner
Nevada Girl	http://en.wikipedia.org/wiki/Nevada_Girl
Neve Campbell	http://en.wikipedia.org/wiki/Neve_Campbell
Nevill F. Mott	http://en.wikipedia.org/wiki/Nevill_F._Mott
Neville Brand	http://en.wikipedia.org/wiki/Neville_Brand
Neville Chamberlain	http://en.wikipedia.org/wiki/Neville_Chamberlain
Newt Gingrich	http://en.wikipedia.org/wiki/Newt_Gingrich
Newt Gingrich	http://en.wikipedia.org/wiki/Newt_Gingrich
Newton D. Baker	http://en.wikipedia.org/wiki/Newton_D._Baker
Nexhat Daci	http://en.wikipedia.org/wiki/Nexhat_Daci
Ngaio Marsh	http://en.wikipedia.org/wiki/Ngaio_Marsh
Nguyen Van Thieu	http://en.wikipedia.org/wiki/Nguyen_Van_Thieu
Nia Griffith	http://en.wikipedia.org/wiki/Nia_Griffith
Nia Long	http://en.wikipedia.org/wiki/Nia_Long
Nia Peeples	http://en.wikipedia.org/wiki/Nia_Peeples
Nia Vardalos	http://en.wikipedia.org/wiki/Nia_Vardalos
Nicanor Duarte	http://en.wikipedia.org/wiki/Nicanor_Duarte
Nicanor Duarte Frutos	http://en.wikipedia.org/wiki/Nicanor_Duarte_Frutos
Niccol� Machiavelli	http://en.wikipedia.org/wiki/Niccol%F2_Machiavelli
Niccol� Niccoli	http://en.wikipedia.org/wiki/Niccol%F2_Niccoli
Niccolo Paganini	http://en.wikipedia.org/wiki/Niccolo_Paganini
Niccol� Tartaglia	http://en.wikipedia.org/wiki/Niccol%F2_Tartaglia
Nicephorus Callistus Xanthopoulos	http://en.wikipedia.org/wiki/Nicephorus_Callistus_Xanthopoulos
Nicephorus I	http://en.wikipedia.org/wiki/Nicephorus_I
Nicephorus II Phocas	http://en.wikipedia.org/wiki/Nicephorus_II_Phocas
Nicephorus III Botaneiates	http://en.wikipedia.org/wiki/Nicephorus_III_Botaneiates
Nicephorus Patriarcha	http://en.wikipedia.org/wiki/Nicephorus_Patriarcha
Nichelle Nichols	http://en.wikipedia.org/wiki/Nichelle_Nichols
Nicholas Amhurst	http://en.wikipedia.org/wiki/Nicholas_Amhurst
Nicholas Biddle	http://en.wikipedia.org/wiki/Nicholas_Biddle_(banker)
Nicholas Brendon	http://en.wikipedia.org/wiki/Nicholas_Brendon
Nicholas Brown	http://en.wikipedia.org/wiki/Nick_Brown
Nicholas Claude Fabri de Peiresc	http://en.wikipedia.org/wiki/Nicolas-Claude_Fabri_de_Peiresc
Nicholas D. Chabraja	http://en.wikipedia.org/wiki/Nicholas_D._Chabraja
Nicholas D. Kristof	http://en.wikipedia.org/wiki/Nicholas_D._Kristof
Nicholas F. Brady	http://en.wikipedia.org/wiki/Nicholas_F._Brady
Nicholas Grimald	http://en.wikipedia.org/wiki/Nicholas_Grimald
Nicholas Hawksmoor	http://en.wikipedia.org/wiki/Nicholas_Hawksmoor
Nicholas Liverpool	http://en.wikipedia.org/wiki/Nicholas_Liverpool
Nicholas Longworth	http://en.wikipedia.org/wiki/Nicholas_Longworth
Nicholas Mavroules	http://en.wikipedia.org/wiki/Nicholas_Mavroules
Nicholas Murray Butler	http://en.wikipedia.org/wiki/Nicholas_Murray_Butler
Nicholas Negroponte	http://en.wikipedia.org/wiki/Nicholas_Negroponte
Nicholas Pileggi	http://en.wikipedia.org/wiki/Nicholas_Pileggi
Nicholas Ray	http://en.wikipedia.org/wiki/Nicholas_Ray
Nicholas Ridley	http://en.wikipedia.org/wiki/Nicholas_Ridley_(martyr)
Nicholas Rowe	http://en.wikipedia.org/wiki/Nicholas_Rowe_(writer)
Nicholas Soames	http://en.wikipedia.org/wiki/Nicholas_Soames
Nicholas Stone	http://en.wikipedia.org/wiki/Nicholas_Stone
Nicholas Turturro	http://en.wikipedia.org/wiki/Nicholas_Turturro
Nick Adams	http://en.wikipedia.org/wiki/Nick_Adams_(actor)
Nick Berg	http://en.wikipedia.org/wiki/Nick_Berg
Nick Boles	http://en.wikipedia.org/wiki/Nick_Boles
Nick Cannon	http://en.wikipedia.org/wiki/Nick_Cannon
Nick Carter	http://en.wikipedia.org/wiki/Nick_Carter_(musician)
Nick Cassavetes	http://en.wikipedia.org/wiki/Nick_Cassavetes
Nick Cave	http://en.wikipedia.org/wiki/Nick_Cave
Nick Clegg	http://en.wikipedia.org/wiki/Nick_Clegg
Nick de Bois	http://en.wikipedia.org/wiki/Nick_de_Bois
Nick Drake	http://en.wikipedia.org/wiki/Nick_Drake
Nick Faldo	http://en.wikipedia.org/wiki/Nick_Faldo
Nick Gibb	http://en.wikipedia.org/wiki/Nick_Gibb
Nick Harvey	http://en.wikipedia.org/wiki/Nick_Harvey
Nick Herbert	http://en.wikipedia.org/wiki/Nick_Herbert
Nick Hornby	http://en.wikipedia.org/wiki/Nick_Hornby
Nick Hurd	http://en.wikipedia.org/wiki/Nick_Hurd
Nick J. Rahall II	http://en.wikipedia.org/wiki/Nick_J._Rahall_II
Nick Lachey	http://en.wikipedia.org/wiki/Nick_Lachey
Nick Lampson	http://en.wikipedia.org/wiki/Nick_Lampson
Nick Lowe	http://en.wikipedia.org/wiki/Nick_Lowe
Nick Mancuso	http://en.wikipedia.org/wiki/Nick_Mancuso
Nick Mason	http://en.wikipedia.org/wiki/Nick_Mason
Nick Nolte	http://en.wikipedia.org/wiki/Nick_Nolte
Nick Oliveri	http://en.wikipedia.org/wiki/Nick_Oliveri
Nick Park	http://en.wikipedia.org/wiki/Nick_Park
Nick Rahall	http://en.wikipedia.org/wiki/Nick_Rahall
Nick Raynsford	http://en.wikipedia.org/wiki/Nick_Raynsford
Nick Rhodes	http://en.wikipedia.org/wiki/Nick_Rhodes
Nick Smith	http://en.wikipedia.org/wiki/Nick_Smith_(U.S._politician)
Nick Smith	http://en.wikipedia.org/wiki/Nick_Smith_(British_politician)
Nick Stahl	http://en.wikipedia.org/wiki/Nick_Stahl
Nick Valensi	http://en.wikipedia.org/wiki/Nick_Valensi
Nick Zano	http://en.wikipedia.org/wiki/Nick_Zano
Nickolas Ashford	http://en.wikipedia.org/wiki/Nickolas_Ashford
Nicky Hilton	http://en.wikipedia.org/wiki/Nicky_Hilton
Nicky Morgan	http://en.wikipedia.org/wiki/Nicky_Morgan_(politician)
Nicol Williamson	http://en.wikipedia.org/wiki/Nicol_Williamson
Nicola Blackwood	http://en.wikipedia.org/wiki/Nicola_Blackwood
Nicola Pisano	http://en.wikipedia.org/wiki/Nicola_Pisano
Nicolaas Bloembergen	http://en.wikipedia.org/wiki/Nicolaas_Bloembergen
Nicolae Ceausescu	http://en.wikipedia.org/wiki/Nicolae_Ceausescu
Nicolas Boileau	http://en.wikipedia.org/wiki/Nicolas_Boileau
Nicolas Cage	http://en.wikipedia.org/wiki/Nicolas_Cage
Nicolas Desmarest	http://en.wikipedia.org/wiki/Nicolas_Desmarest
Nicolas Godin	http://en.wikipedia.org/wiki/Nicolas_Godin
Nicolas Jenson	http://en.wikipedia.org/wiki/Nicolas_Jenson
Nicolas Louis de Lacaille	http://en.wikipedia.org/wiki/Nicolas_Louis_de_Lacaille
Nicolas Malebranche	http://en.wikipedia.org/wiki/Nicolas_Malebranche
Nicolas Poussin	http://en.wikipedia.org/wiki/Nicolas_Poussin
Nicolas Roeg	http://en.wikipedia.org/wiki/Nicolas_Roeg
Nicolas Sarkozy	http://en.wikipedia.org/wiki/Nicolas_Sarkozy
Nicolas-Charles Oudinot	http://en.wikipedia.org/wiki/Nicolas_Oudinot
Nicolas-Louis Vauquelin	http://en.wikipedia.org/wiki/Nicolas-Louis_Vauquelin
Nicolaus Copernicus	http://en.wikipedia.org/wiki/Nicolaus_Copernicus
Nicolaus Steno	http://en.wikipedia.org/wiki/Nicolaus_Steno
Nicole Appleton	http://en.wikipedia.org/wiki/Nicole_Appleton
Nicole Ari Parker	http://en.wikipedia.org/wiki/Nicole_Ari_Parker
Nicole Brown Simpson	http://en.wikipedia.org/wiki/Nicole_Brown_Simpson
Nicole DeHuff	http://en.wikipedia.org/wiki/Nicole_DeHuff
Nicole Eggert	http://en.wikipedia.org/wiki/Nicole_Eggert
Nicole Holofcener	http://en.wikipedia.org/wiki/Nicole_Holofcener
Nicole Kidman	http://en.wikipedia.org/wiki/Nicole_Kidman
Nicole Richie	http://en.wikipedia.org/wiki/Nicole_Richie
Nicole Scherzinger	http://en.wikipedia.org/wiki/Nicole_Scherzinger
Nicole Sullivan	http://en.wikipedia.org/wiki/Nicole_Sullivan
Nicolette Sheridan	http://en.wikipedia.org/wiki/Nicolette_Sheridan
Niecy Nash	http://en.wikipedia.org/wiki/Niecy_Nash
Niels Bohr	http://en.wikipedia.org/wiki/Niels_Bohr
Niels Henrik Abel	http://en.wikipedia.org/wiki/Niels_Henrik_Abel
Niels Ryberg Finsen	http://en.wikipedia.org/wiki/Niels_Ryberg_Finsen
Nigel Adams	http://en.wikipedia.org/wiki/Nigel_Adams
Nigel Bruce	http://en.wikipedia.org/wiki/Nigel_Bruce
Nigel Dennis	http://en.wikipedia.org/wiki/Nigel_Dennis
Nigel Dodds	http://en.wikipedia.org/wiki/Nigel_Dodds
Nigel Evans	http://en.wikipedia.org/wiki/Nigel_Evans
Nigel Godrich	http://en.wikipedia.org/wiki/Nigel_Godrich
Nigel Hawthorne	http://en.wikipedia.org/wiki/Nigel_Hawthorne
Nigel Kennedy	http://en.wikipedia.org/wiki/Nigel_Kennedy
Nigel Mills	http://en.wikipedia.org/wiki/Nigel_Mills
Nigella Lawson	http://en.wikipedia.org/wiki/Nigella_Lawson
Nik Kershaw	http://en.wikipedia.org/wiki/Nik_Kershaw
Niki Sullivan	http://en.wikipedia.org/wiki/Niki_Sullivan
Niki Taylor	http://en.wikipedia.org/wiki/Niki_Taylor
Niki Tsongas	http://en.wikipedia.org/wiki/Niki_Tsongas
Nikita Khrushchev	http://en.wikipedia.org/wiki/Nikita_Khrushchev
Nikki Amuka-Bird	http://en.wikipedia.org/wiki/Nikki_Amuka-Bird
Nikki Cox	http://en.wikipedia.org/wiki/Nikki_Cox
Nikki Fritz	http://en.wikipedia.org/wiki/Nikki_Fritz
Nikki Giovanni	http://en.wikipedia.org/wiki/Nikki_Giovanni
Nikki Reed	http://en.wikipedia.org/wiki/Nikki_Reed
Nikki Sixx	http://en.wikipedia.org/wiki/Nikki_Sixx
Niklaus Wirth	http://en.wikipedia.org/wiki/Niklaus_Wirth
Niko Lozancic	http://en.wikipedia.org/wiki/Niko_Lozancic
Nikola Gruevski	http://en.wikipedia.org/wiki/Nikola_Gruevski
Nikola Tesla	http://en.wikipedia.org/wiki/Nikola_Tesla
Nikolaas Tinbergen	http://en.wikipedia.org/wiki/Nikolaas_Tinbergen
Nikolai Cherkasov	http://en.wikipedia.org/wiki/Nikolai_Cherkasov
Nikolai Dzhurmongaliev	http://en.wikipedia.org/wiki/Nikolai_Dzhurmongaliev
Nikolai Fraiture	http://en.wikipedia.org/wiki/Nikolai_Fraiture
Nikolai Gogol	http://en.wikipedia.org/wiki/Nikolai_Gogol
Nikolai Novikov	http://en.wikipedia.org/wiki/Nikolai_Novikov
Nikolai Podgorny	http://en.wikipedia.org/wiki/Nikolai_Podgorny
Nikolai Rimsky-Korsakov	http://en.wikipedia.org/wiki/Nikolai_Rimsky-Korsakov
Nikolai Ryzhkov	http://en.wikipedia.org/wiki/Nikolai_Ryzhkov
Nikolai Tikhonov	http://en.wikipedia.org/wiki/Nikolai_Tikhonov
Nikolai Yazykov	http://en.wikipedia.org/wiki/Nikolai_Yazykov
Nikolaus von Amsdorf	http://en.wikipedia.org/wiki/Nikolaus_von_Amsdorf
Nikolay G. Basov	http://en.wikipedia.org/wiki/Nikolay_Basov
Nikolay Semyonov	http://en.wikipedia.org/wiki/Nikolay_Semyonov
Nikoloz Gilauri	http://en.wikipedia.org/wiki/Nikoloz_Gilauri
Nikos Kazantzakis	http://en.wikipedia.org/wiki/Nikos_Kazantzakis
Nile Rodgers	http://en.wikipedia.org/wiki/Nile_Rodgers
Nils Asther	http://en.wikipedia.org/wiki/Nils_Asther
Nils Frykdahl	http://en.wikipedia.org/wiki/Nils_Frykdahl
Nils Lofgren	http://en.wikipedia.org/wiki/Nils_Lofgren
Nina Alisova	http://en.wikipedia.org/wiki/Nina_Alisova
Nina Bawden	http://en.wikipedia.org/wiki/Nina_Bawden
Nina Blackwood	http://en.wikipedia.org/wiki/Nina_Blackwood
Nina Foch	http://en.wikipedia.org/wiki/Nina_Foch
Nina Hagen	http://en.wikipedia.org/wiki/Nina_Hagen
Nina Munk	http://en.wikipedia.org/wiki/Nina_Munk
Nina Simone	http://en.wikipedia.org/wiki/Nina_Simone
Nina Totenberg	http://en.wikipedia.org/wiki/Nina_Totenberg
Nino Rota	http://en.wikipedia.org/wiki/Nino_Rota
Nipsey Russell	http://en.wikipedia.org/wiki/Nipsey_Russell
Nita Lowey	http://en.wikipedia.org/wiki/Nita_Lowey
Nivek Ogre	http://en.wikipedia.org/wiki/Nivek_Ogre
NO I.D.	http://en.wikipedia.org/wiki/NO_I.D.
Noah Adams	http://en.wikipedia.org/wiki/Noah_Adams
Noah Beery, Jr.	http://en.wikipedia.org/wiki/Noah_Beery%2C_Jr.
Noah Beery, Sr.	http://en.wikipedia.org/wiki/Noah_Beery%2C_Sr.
Noah Hathaway	http://en.wikipedia.org/wiki/Noah_Hathaway
Noah Kadner	http://en.wikipedia.org/wiki/Noah_Kadner
Noah Taylor	http://en.wikipedia.org/wiki/Noah_Taylor
Noah Webster	http://en.wikipedia.org/wiki/Noah_Webster
Noah Wyle	http://en.wikipedia.org/wiki/Noah_Wyle
Noam Chomsky	http://en.wikipedia.org/wiki/Noam_Chomsky
Noble Willingham	http://en.wikipedia.org/wiki/Noble_Willingham
Nobuo Uematsu	http://en.wikipedia.org/wiki/Nobuo_Uematsu
Noel Coward	http://en.wikipedia.org/wiki/Noel_Coward
No�l Forgeard	http://en.wikipedia.org/wiki/No%EBl_Forgeard
Noel Gallagher	http://en.wikipedia.org/wiki/Noel_Gallagher
Noel Redding	http://en.wikipedia.org/wiki/Noel_Redding
Noelle Bush	http://en.wikipedia.org/wiki/Noelle_Bush
Nolan Bushnell	http://en.wikipedia.org/wiki/Nolan_Bushnell
Nolan Ryan	http://en.wikipedia.org/wiki/Nolan_Ryan
Nomar Garciaparra	http://en.wikipedia.org/wiki/Nomar_Garciaparra
Nona Gaye	http://en.wikipedia.org/wiki/Nona_Gaye
Nona Hendryx	http://en.wikipedia.org/wiki/Nona_Hendryx
Nong Duc Manh	http://en.wikipedia.org/wiki/Nong_Duc_Manh
Nora Dunn	http://en.wikipedia.org/wiki/Nora_Dunn
Nora Ephron	http://en.wikipedia.org/wiki/Nora_Ephron
Norah Jones	http://en.wikipedia.org/wiki/Norah_Jones
Norbert Wiener	http://en.wikipedia.org/wiki/Norbert_Wiener
Norm Abram	http://en.wikipedia.org/wiki/Norm_Abram
Norm Coleman	http://en.wikipedia.org/wiki/Norm_Coleman
Norm Crosby	http://en.wikipedia.org/wiki/Norm_Crosby
Norm Dicks	http://en.wikipedia.org/wiki/Norm_Dicks
Norm MacDonald	http://en.wikipedia.org/wiki/Norm_MacDonald_(comedian)
Norm Mineta	http://en.wikipedia.org/wiki/Norm_Mineta
Norma Khouri	http://en.wikipedia.org/wiki/Norma_Khouri
Norma McCorvey	http://en.wikipedia.org/wiki/Norma_McCorvey
Norma Shearer	http://en.wikipedia.org/wiki/Norma_Shearer
Norman Angell	http://en.wikipedia.org/wiki/Norman_Angell
Norman Augustine	http://en.wikipedia.org/wiki/Norman_Augustine
Norman Baker	http://en.wikipedia.org/wiki/Norman_Baker
Norman Borlaug	http://en.wikipedia.org/wiki/Norman_Borlaug
Norman Campbell	http://en.wikipedia.org/wiki/Norman_Campbell
Norman Cousins	http://en.wikipedia.org/wiki/Norman_Cousins
Norman D. Dicks	http://en.wikipedia.org/wiki/Norman_D._Dicks
Norman D. Shumway	http://en.wikipedia.org/wiki/Norman_D._Shumway
Norman Dello Joio	http://en.wikipedia.org/wiki/Norman_Dello_Joio
Norman F. Lent	http://en.wikipedia.org/wiki/Norman_F._Lent
Norman F. Ramsey	http://en.wikipedia.org/wiki/Norman_F._Ramsey
Norman Fell	http://en.wikipedia.org/wiki/Norman_Fell
Norman Foster	http://en.wikipedia.org/wiki/Norman_Foster_(architect)
Norman Haworth	http://en.wikipedia.org/wiki/Norman_Haworth
Norman Jewison	http://en.wikipedia.org/wiki/Norman_Jewison
Norman Lamb	http://en.wikipedia.org/wiki/Norman_Lamb
Norman Lear	http://en.wikipedia.org/wiki/Norman_Lear
Norman Lloyd	http://en.wikipedia.org/wiki/Norman_Lloyd
Norman Mailer	http://en.wikipedia.org/wiki/Norman_Mailer
Norman Ornstein	http://en.wikipedia.org/wiki/Norman_Ornstein
Norman Parker	http://en.wikipedia.org/wiki/Norman_Parker
Norman Podhoretz	http://en.wikipedia.org/wiki/Norman_Podhoretz
Norman Reedus	http://en.wikipedia.org/wiki/Norman_Reedus
Norman Rockwell	http://en.wikipedia.org/wiki/Norman_Rockwell
Norman Rush	http://en.wikipedia.org/wiki/Norman_Rush
Norman Schwarzkopf	http://en.wikipedia.org/wiki/Norman_Schwarzkopf
Norman Sisisky	http://en.wikipedia.org/wiki/Norman_Sisisky
Norman Spinrad	http://en.wikipedia.org/wiki/Norman_Spinrad
Norman Taurog	http://en.wikipedia.org/wiki/Norman_Taurog
Norman Tokar	http://en.wikipedia.org/wiki/Norman_Tokar
Norman Vincent Peale	http://en.wikipedia.org/wiki/Norman_Vincent_Peale
Norman Wisdom	http://en.wikipedia.org/wiki/Norman_Wisdom
Norman Y. Mineta	http://en.wikipedia.org/wiki/Norman_Y._Mineta
Norman Z. McLeod	http://en.wikipedia.org/wiki/Norman_Z._McLeod
Norodom Sihanouk	http://en.wikipedia.org/wiki/Norodom_Sihanouk
Norris Church Mailer	http://en.wikipedia.org/wiki/Norris_Church_Mailer
Norris McWhirter	http://en.wikipedia.org/wiki/Norris_McWhirter
Norris Poulson	http://en.wikipedia.org/wiki/Norris_Poulson
Northrop Frye	http://en.wikipedia.org/wiki/Northrop_Frye
Norton Juster	http://en.wikipedia.org/wiki/Norton_Juster
Norton Schwartz	http://en.wikipedia.org/wiki/Norton_Schwartz
Norton Simon	http://en.wikipedia.org/wiki/Norton_Simon
Notorious B.I.G.	http://en.wikipedia.org/wiki/Notorious_B.I.G.
Nouri al-Maliki	http://en.wikipedia.org/wiki/Nouri_al-Maliki
Nunnally Johnson	http://en.wikipedia.org/wiki/Nunnally_Johnson
Nuno Bettencourt	http://en.wikipedia.org/wiki/Nuno_Bettencourt
Nur Muhammad Taraki	http://en.wikipedia.org/wiki/Nur_Muhammad_Taraki
Nuri al-Maliki	http://en.wikipedia.org/wiki/Nuri_al-Maliki
Nursultan Nazarbayev	http://en.wikipedia.org/wiki/Nursultan_Nazarbayev
Nuruddin Farah	http://en.wikipedia.org/wiki/Nuruddin_Farah
Nusrat Fateh Ali Khan	http://en.wikipedia.org/wiki/Nusrat_Fateh_Ali_Khan
Nydia Vel�zquez	http://en.wikipedia.org/wiki/Nydia_Vel%E1zquez
Nyree Dawn Porter	http://en.wikipedia.org/wiki/Nyree_Dawn_Porter
O. E. R�lvaag	http://en.wikipedia.org/wiki/Ole_Edvart_R%C3%B8lvaag
O. Henry	http://en.wikipedia.org/wiki/O._Henry
O. J. Simpson	http://en.wikipedia.org/wiki/O._J._Simpson
Obba Babatund�	http://en.wikipedia.org/wiki/Obba_Babatund%E9
Obie Trice	http://en.wikipedia.org/wiki/Obie_Trice
Octavia Butler	http://en.wikipedia.org/wiki/Octavia_Butler
Octavio Paz	http://en.wikipedia.org/wiki/Octavio_Paz
Odd Hassel	http://en.wikipedia.org/wiki/Odd_Hassel
Oded Fehr	http://en.wikipedia.org/wiki/Oded_Fehr
Odilon Redon	http://en.wikipedia.org/wiki/Odilon_Redon
Odo of Bayeux	http://en.wikipedia.org/wiki/Odo_of_Bayeux
Ogden Nash	http://en.wikipedia.org/wiki/Ogden_Nash
Ogi Ogas	http://en.wikipedia.org/wiki/Ogi_Ogas
Oksana Baiul	http://en.wikipedia.org/wiki/Oksana_Baiul
Ol' Dirty Bastard	http://en.wikipedia.org/wiki/Ol%27_Dirty_Bastard
Olaf I Tryggvason	http://en.wikipedia.org/wiki/Olaf_I_Tryggvason
Olaf II Haraldsson	http://en.wikipedia.org/wiki/Olaf_II_Haraldsson
�lafur Ragnar Gr�msson	http://en.wikipedia.org/wiki/%D3lafur_Ragnar_Gr%EDmsson
Olaus Magnus	http://en.wikipedia.org/wiki/Olaus_Magnus
Oleg Cassini	http://en.wikipedia.org/wiki/Oleg_Cassini
Olene Walker	http://en.wikipedia.org/wiki/Olene_Walker
Olga Korbut	http://en.wikipedia.org/wiki/Olga_Korbut
Olive Carey	http://en.wikipedia.org/wiki/Olive_Carey
Olive Schreiner	http://en.wikipedia.org/wiki/Olive_Schreiner
Oliver Colvile	http://en.wikipedia.org/wiki/Oliver_Colvile
Oliver Cromwell	http://en.wikipedia.org/wiki/Oliver_Cromwell
Oliver Goldsmith	http://en.wikipedia.org/wiki/Oliver_Goldsmith
Oliver Hardy	http://en.wikipedia.org/wiki/Oliver_Hardy
Oliver Hazard Perry	http://en.wikipedia.org/wiki/Oliver_Hazard_Perry
Oliver Heald	http://en.wikipedia.org/wiki/Oliver_Heald
Oliver Herford	http://en.wikipedia.org/wiki/Oliver_Herford
Oliver Hudson	http://en.wikipedia.org/wiki/Oliver_Hudson
Oliver James	http://en.wikipedia.org/wiki/Oliver_James_(entertainer)
Oliver La Farge	http://en.wikipedia.org/wiki/Oliver_La_Farge
Oliver Letwin	http://en.wikipedia.org/wiki/Oliver_Letwin
Oliver North	http://en.wikipedia.org/wiki/Oliver_North
Oliver O. Howard	http://en.wikipedia.org/wiki/Oliver_O._Howard
Oliver Perry Morton	http://en.wikipedia.org/wiki/Oliver_Perry_Morton
Oliver Platt	http://en.wikipedia.org/wiki/Oliver_Platt
Oliver Reed	http://en.wikipedia.org/wiki/Oliver_Reed
Oliver Stone	http://en.wikipedia.org/wiki/Oliver_Stone
Oliver Tambo	http://en.wikipedia.org/wiki/Oliver_Tambo
Oliver Wendell Holmes	http://en.wikipedia.org/wiki/Oliver_Wendell_Holmes
Oliver Wendell Holmes, Jr.	http://en.wikipedia.org/wiki/Oliver_Wendell_Holmes%2C_Jr.
Olivia d'Abo	http://en.wikipedia.org/wiki/Olivia_d%27Abo
Olivia de Havilland	http://en.wikipedia.org/wiki/Olivia_de_Havilland
Olivia de Havilland	http://en.wikipedia.org/wiki/Olivia_de_Havilland
Olivia Goldsmith	http://en.wikipedia.org/wiki/Olivia_Goldsmith
Olivia Hussey	http://en.wikipedia.org/wiki/Olivia_Hussey
Olivia Newton-John	http://en.wikipedia.org/wiki/Olivia_Newton-John
Olivia Wilde	http://en.wikipedia.org/wiki/Olivia_Wilde
Olivier Martinez	http://en.wikipedia.org/wiki/Olivier_Martinez
Olivier Messiaen	http://en.wikipedia.org/wiki/Olivier_Messiaen
Olle Adolphson	http://en.wikipedia.org/wiki/Olle_Adolphson
Olof Palme	http://en.wikipedia.org/wiki/Olof_Palme
Olusegun Obasanjo	http://en.wikipedia.org/wiki/Olusegun_Obasanjo
Olusegun Obasanjo	http://en.wikipedia.org/wiki/Olusegun_Obasanjo
Olympia Dukakis	http://en.wikipedia.org/wiki/Olympia_Dukakis
Olympia J. Snowe	http://en.wikipedia.org/wiki/Olympia_J._Snowe
Olympia Snowe	http://en.wikipedia.org/wiki/Olympia_Snowe
Omar Abdel-Rahman	http://en.wikipedia.org/wiki/Omar_Abdel-Rahman
Omar Abdirashid Ali Sharmarke	http://en.wikipedia.org/wiki/Omar_Abdirashid_Ali_Sharmarke
Omar al-Bashir	http://en.wikipedia.org/wiki/Omar_al-Bashir
Omar Al-Qattan	http://en.wikipedia.org/wiki/Omar_Al-Qattan
Omar Bongo	http://en.wikipedia.org/wiki/Omar_Bongo
Omar Bradley	http://en.wikipedia.org/wiki/Omar_Bradley
Omar Epps	http://en.wikipedia.org/wiki/Omar_Epps
Omar Gooding	http://en.wikipedia.org/wiki/Omar_Gooding
Omar Hasan Ahmad al-Bashir	http://en.wikipedia.org/wiki/Omar_Hasan_Ahmad_al-Bashir
Omar Khayyam	http://en.wikipedia.org/wiki/Omar_Khayyam
Omar Sharif	http://en.wikipedia.org/wiki/Omar_Sharif
Omar Torrijos	http://en.wikipedia.org/wiki/Omar_Torrijos
Omri Katz	http://en.wikipedia.org/wiki/Omri_Katz
Opie Read	http://en.wikipedia.org/wiki/Opie_Read
Oprah Winfrey	http://en.wikipedia.org/wiki/Oprah_Winfrey
Oqil Oqilov	http://en.wikipedia.org/wiki/Oqil_Oqilov
Oral Roberts	http://en.wikipedia.org/wiki/Oral_Roberts
Orazio Gentileschi	http://en.wikipedia.org/wiki/Orazio_Gentileschi
Orel Hershiser	http://en.wikipedia.org/wiki/Orel_Hershiser
Orhan I	http://en.wikipedia.org/wiki/Orhan_I
Orhan Pamuk	http://en.wikipedia.org/wiki/Orhan_Pamuk
Orin C. Smith	http://en.wikipedia.org/wiki/Orin_C._Smith
Orkut Buyukkokten	http://en.wikipedia.org/wiki/Orkut_Buyukkokten
Orlando Bloom	http://en.wikipedia.org/wiki/Orlando_Bloom
Orlando Brown	http://en.wikipedia.org/wiki/Orlando_Brown
Orlando di Lasso	http://en.wikipedia.org/wiki/Orlando_di_Lasso
Orlando Gibbons	http://en.wikipedia.org/wiki/Orlando_Gibbons
Orlando Jones	http://en.wikipedia.org/wiki/Orlando_Jones
Ornette Coleman	http://en.wikipedia.org/wiki/Ornette_Coleman
Orrin G. Hatch	http://en.wikipedia.org/wiki/Orrin_G._Hatch
Orrin Hatch	http://en.wikipedia.org/wiki/Orrin_Hatch
Orson Bean	http://en.wikipedia.org/wiki/Orson_Bean
Orson Scott Card	http://en.wikipedia.org/wiki/Orson_Scott_Card
Orson Welles	http://en.wikipedia.org/wiki/Orson_Welles
Orville Wright	http://en.wikipedia.org/wiki/Orville_Wright
Osama bin Laden	http://en.wikipedia.org/wiki/Osama_bin_Laden
Osamu Akimoto	http://en.wikipedia.org/wiki/Osamu_Akimoto
�scar Arias	http://en.wikipedia.org/wiki/%D3scar_Arias
Oscar Arias Sanchez	http://en.wikipedia.org/wiki/Oscar_Arias_Sanchez
�scar Berger	http://en.wikipedia.org/wiki/%D3scar_Berger
Oscar De La Hoya	http://en.wikipedia.org/wiki/Oscar_De_La_Hoya
Oscar de la Renta	http://en.wikipedia.org/wiki/Oscar_de_la_Renta
Oscar Hammerstein	http://en.wikipedia.org/wiki/Oscar_Hammerstein_II
Oscar Handlin	http://en.wikipedia.org/wiki/Oscar_Handlin
Oscar Hijuelos	http://en.wikipedia.org/wiki/Oscar_Hijuelos
Oscar I	http://en.wikipedia.org/wiki/Oscar_I
Oscar II	http://en.wikipedia.org/wiki/Oscar_II_of_Sweden
Oscar L. Chapman	http://en.wikipedia.org/wiki/Oscar_L._Chapman
Oscar Mayer	http://en.wikipedia.org/wiki/Oscar_F._Mayer
Oscar Niemeyer	http://en.wikipedia.org/wiki/Oscar_Niemeyer
Oscar Robertson	http://en.wikipedia.org/wiki/Oscar_Robertson
Oscar Temaru	http://en.wikipedia.org/wiki/Oscar_Temaru
Oscar Wilde	http://en.wikipedia.org/wiki/Oscar_Wilde
Osip Mandelshtam	http://en.wikipedia.org/wiki/Osip_Mandelshtam
Oskar Kokoschka	http://en.wikipedia.org/wiki/Oskar_Kokoschka
Oskar Schindler	http://en.wikipedia.org/wiki/Oskar_Schindler
Osman I	http://en.wikipedia.org/wiki/Osman_I
Ossie Davis	http://en.wikipedia.org/wiki/Ossie_Davis
Oswald Mosley	http://en.wikipedia.org/wiki/Oswald_Mosley
Oswald Myconius	http://en.wikipedia.org/wiki/Oswald_Myconius
Oswald Spengler	http://en.wikipedia.org/wiki/Oswald_Spengler
Otis Blackwell	http://en.wikipedia.org/wiki/Otis_Blackwell
Otis Chandler	http://en.wikipedia.org/wiki/Otis_Chandler
Otis Redding	http://en.wikipedia.org/wiki/Otis_Redding
Otis Williams	http://en.wikipedia.org/wiki/Otis_Williams
Otmar Hasler	http://en.wikipedia.org/wiki/Otmar_Hasler
Otto Diels	http://en.wikipedia.org/wiki/Otto_Diels
Otto Dix	http://en.wikipedia.org/wiki/Otto_Dix
Otto Hahn	http://en.wikipedia.org/wiki/Otto_Hahn
Otto I	http://en.wikipedia.org/wiki/Otto_I
Otto II	http://en.wikipedia.org/wiki/Otto_II
Otto III	http://en.wikipedia.org/wiki/Otto_III
Otto IV	http://en.wikipedia.org/wiki/Otto_IV
Otto Kahn	http://en.wikipedia.org/wiki/Otto_Kahn
Otto Klemperer	http://en.wikipedia.org/wiki/Otto_Klemperer
Otto Kruger	http://en.wikipedia.org/wiki/Otto_Kruger
Otto Ludwig	http://en.wikipedia.org/wiki/Otto_Ludwig_(writer)
Otto Neurath	http://en.wikipedia.org/wiki/Otto_Neurath
Otto of Freising	http://en.wikipedia.org/wiki/Otto_of_Freising
Otto Preminger	http://en.wikipedia.org/wiki/Otto_Preminger
Otto Robert Frisch	http://en.wikipedia.org/wiki/Otto_Robert_Frisch
Otto Schily	http://en.wikipedia.org/wiki/Otto_Schily
Otto Skorzeny	http://en.wikipedia.org/wiki/Otto_Skorzeny
Otto Stern	http://en.wikipedia.org/wiki/Otto_Stern
Otto von Bismarck	http://en.wikipedia.org/wiki/Otto_von_Bismarck
Otto Wallach	http://en.wikipedia.org/wiki/Otto_Wallach
Otto Wilhelm Struve	http://en.wikipedia.org/wiki/Otto_Wilhelm_Struve
Ottorino Respighi	http://en.wikipedia.org/wiki/Ottorino_Respighi
Ousmane Issoufi Ma�ga	http://en.wikipedia.org/wiki/Ousmane_Issoufi_Ma%EFga
Ove Arup	http://en.wikipedia.org/wiki/Ove_Arup
Owen Arthur	http://en.wikipedia.org/wiki/Owen_Arthur
Owen Chamberlain	http://en.wikipedia.org/wiki/Owen_Chamberlain
Owen Glendower	http://en.wikipedia.org/wiki/Owen_Glendower
Owen Hart	http://en.wikipedia.org/wiki/Owen_Hart
Owen Paterson	http://en.wikipedia.org/wiki/Owen_Paterson
Owen Smith	http://en.wikipedia.org/wiki/Owen_Smith
Owen Willans Richardson	http://en.wikipedia.org/wiki/Owen_Willans_Richardson
Owen Wilson	http://en.wikipedia.org/wiki/Owen_Wilson
Owen Wister	http://en.wikipedia.org/wiki/Owen_Wister
Owsley Stanley	http://en.wikipedia.org/wiki/Owsley_Stanley
Ozzie Nelson	http://en.wikipedia.org/wiki/Ozzie_Nelson
Ozzie Smith	http://en.wikipedia.org/wiki/Ozzie_Smith
Ozzy Osbourne	http://en.wikipedia.org/wiki/Ozzy_Osbourne
P. D. James	http://en.wikipedia.org/wiki/P._D._James
P. G. Wodehouse	http://en.wikipedia.org/wiki/P._G._Wodehouse
P. J. Harvey	http://en.wikipedia.org/wiki/P._J._Harvey
P. J. O'Rourke	http://en.wikipedia.org/wiki/P._J._O%27Rourke
P. P. Arnold	http://en.wikipedia.org/wiki/P._P._Arnold
P. T. Barnum	http://en.wikipedia.org/wiki/P._T._Barnum
P. W. Botha	http://en.wikipedia.org/wiki/P._W._Botha
P.J. Patterson	http://en.wikipedia.org/wiki/P.J._Patterson
Pablo Casals	http://en.wikipedia.org/wiki/Pablo_Casals
Pablo de C�spedes	http://en.wikipedia.org/wiki/Pablo_de_C%E9spedes
Pablo Escobar	http://en.wikipedia.org/wiki/Pablo_Escobar
Pablo Neruda	http://en.wikipedia.org/wiki/Pablo_Neruda
Pablo Picasso	http://en.wikipedia.org/wiki/Pablo_Picasso
Paddy Ashdown	http://en.wikipedia.org/wiki/Paddy_Ashdown
Paddy Chayefsky	http://en.wikipedia.org/wiki/Paddy_Chayefsky
Padraic Colum	http://en.wikipedia.org/wiki/Padraic_Colum
Page McConnell	http://en.wikipedia.org/wiki/Page_McConnell
Paige Davis	http://en.wikipedia.org/wiki/Paige_Davis
Pak Pong-ju	http://en.wikipedia.org/wiki/Pak_Pong-ju
Pakalitha Mosisili	http://en.wikipedia.org/wiki/Pakalitha_Mosisili
Pam Dawber	http://en.wikipedia.org/wiki/Pam_Dawber
Pam Grier	http://en.wikipedia.org/wiki/Pam_Grier
Pamela Anderson	http://en.wikipedia.org/wiki/Pamela_Anderson
Pamela Anderson Lee	http://en.wikipedia.org/wiki/Pamela_Anderson_Lee
Pamela Harriman	http://en.wikipedia.org/wiki/Pamela_Harriman
Pamela Nash	http://en.wikipedia.org/wiki/Pamela_Nash
Pamela S. Karlan	http://en.wikipedia.org/wiki/Pamela_S._Karlan
Pamela Segall	http://en.wikipedia.org/wiki/Pamela_Segall
Pamela Stephenson	http://en.wikipedia.org/wiki/Pamela_Stephenson
Pamela Sue Martin	http://en.wikipedia.org/wiki/Pamela_Sue_Martin
Pamela Tiffin	http://en.wikipedia.org/wiki/Pamela_Tiffin
Pancho Villa	http://en.wikipedia.org/wiki/Pancho_Villa
Pandeli Majko	http://en.wikipedia.org/wiki/Pandeli_Majko
Pandro S. Berman	http://en.wikipedia.org/wiki/Pandro_S._Berman
Paolo Di Canio	http://en.wikipedia.org/wiki/Paolo_Di_Canio
Paolo Maldini	http://en.wikipedia.org/wiki/Paolo_Maldini
Paolo Paruta	http://en.wikipedia.org/wiki/Paolo_Paruta
Paolo Sarpi	http://en.wikipedia.org/wiki/Paolo_Sarpi
Paolo Uccello	http://en.wikipedia.org/wiki/Paolo_Uccello
Paolo Veronese	http://en.wikipedia.org/wiki/Paolo_Veronese
Papa Wemba	http://en.wikipedia.org/wiki/Papa_Wemba
P�r Lagerkvist	http://en.wikipedia.org/wiki/P%E4r_Lagerkvist
Paramanga Ernest Yonli	http://en.wikipedia.org/wiki/Paramanga_Ernest_Yonli
Paris Bordone	http://en.wikipedia.org/wiki/Paris_Bordone
Paris Hilton	http://en.wikipedia.org/wiki/Paris_Hilton
Paris Latsis	http://en.wikipedia.org/wiki/Paris_Latsis
Park Chung Hee	http://en.wikipedia.org/wiki/Park_Chung_Hee
Parker Griffith	http://en.wikipedia.org/wiki/Parker_Griffith
Parker Posey	http://en.wikipedia.org/wiki/Parker_Posey
Parker Stevenson	http://en.wikipedia.org/wiki/Parker_Stevenson
Parminder Nagra	http://en.wikipedia.org/wiki/Parminder_Nagra
Parren J. Mitchell	http://en.wikipedia.org/wiki/Parren_J._Mitchell
Parveen Babi	http://en.wikipedia.org/wiki/Parveen_Babi
Pascal Yoadimnadji	http://en.wikipedia.org/wiki/Pascal_Yoadimnadji
Pascual Jordan	http://en.wikipedia.org/wiki/Pascual_Jordan
Pasqual Maragall i Mira	http://en.wikipedia.org/wiki/Pasqual_Maragall_i_Mira
Pasquale Paoli	http://en.wikipedia.org/wiki/Pasquale_Paoli
Pat Barker	http://en.wikipedia.org/wiki/Pat_Barker
Pat Benatar	http://en.wikipedia.org/wiki/Pat_Benatar
Pat Boone	http://en.wikipedia.org/wiki/Pat_Boone
Pat Brown	http://en.wikipedia.org/wiki/Pat_Brown
Pat Buchanan	http://en.wikipedia.org/wiki/Pat_Buchanan
Pat Conroy	http://en.wikipedia.org/wiki/Pat_Conroy
Pat Doherty	http://en.wikipedia.org/wiki/Pat_Doherty
Pat Glass	http://en.wikipedia.org/wiki/Pat_Glass
Pat Harrington, Jr.	http://en.wikipedia.org/wiki/Pat_Harrington%2C_Jr.
Pat Hingle	http://en.wikipedia.org/wiki/Pat_Hingle
Pat Mastelotto	http://en.wikipedia.org/wiki/Pat_Mastelotto
Pat McCarran	http://en.wikipedia.org/wiki/Pat_McCarran
Pat McFadden	http://en.wikipedia.org/wiki/Pat_McFadden_(British_politician)
Pat Metheny	http://en.wikipedia.org/wiki/Pat_Metheny
Pat Morita	http://en.wikipedia.org/wiki/Pat_Morita
Pat Nixon	http://en.wikipedia.org/wiki/Pat_Nixon
Pat O'Brien	http://en.wikipedia.org/wiki/Pat_O'Brien_(television)
Pat O'Brien	http://en.wikipedia.org/wiki/Pat_O'Brien_(actor)
Pat Oliphant	http://en.wikipedia.org/wiki/Pat_Oliphant
Pat Priest	http://en.wikipedia.org/wiki/Pat_Priest
Pat Roberts	http://en.wikipedia.org/wiki/Pat_Roberts
Pat Roberts	http://en.wikipedia.org/wiki/Pat_Roberts
Pat Robertson	http://en.wikipedia.org/wiki/Pat_Robertson
Pat Sajak	http://en.wikipedia.org/wiki/Pat_Sajak
Pat Schroeder	http://en.wikipedia.org/wiki/Pat_Schroeder
Pat Smear	http://en.wikipedia.org/wiki/Pat_Smear
Pat Summerall	http://en.wikipedia.org/wiki/Pat_Summerall
Pat Swindall	http://en.wikipedia.org/wiki/Pat_Swindall
Pat Tiberi	http://en.wikipedia.org/wiki/Pat_Tiberi
Pat Tillman	http://en.wikipedia.org/wiki/Pat_Tillman
Pat Toomey	http://en.wikipedia.org/wiki/Pat_Toomey
Pat Travers	http://en.wikipedia.org/wiki/Pat_Travers
Pat Williams	http://en.wikipedia.org/wiki/John_Patrick_Williams
Patric Knowles	http://en.wikipedia.org/wiki/Patric_Knowles
Patrice Lumumba	http://en.wikipedia.org/wiki/Patrice_Lumumba
Patricia Arquette	http://en.wikipedia.org/wiki/Patricia_Arquette
Patricia Clarkson	http://en.wikipedia.org/wiki/Patricia_Clarkson
Patricia Cornwell	http://en.wikipedia.org/wiki/Patricia_Cornwell
Patricia F. Russo	http://en.wikipedia.org/wiki/Patricia_F._Russo
Patricia Ford	http://en.wikipedia.org/wiki/Patricia_Ford
Patricia Heaton	http://en.wikipedia.org/wiki/Patricia_Heaton
Patricia Highsmith	http://en.wikipedia.org/wiki/Patricia_Highsmith
Patricia Ireland	http://en.wikipedia.org/wiki/Patricia_Ireland
Patricia Medina	http://en.wikipedia.org/wiki/Patricia_Medina
Patricia Neal	http://en.wikipedia.org/wiki/Patricia_Neal
Patricia Quinn	http://en.wikipedia.org/wiki/Patricia_Quinn
Patricia Richardson	http://en.wikipedia.org/wiki/Patricia_Richardson
Patricia Roc	http://en.wikipedia.org/wiki/Patricia_Roc
Patricia Routledge	http://en.wikipedia.org/wiki/Patricia_Routledge
Patricia Schroeder	http://en.wikipedia.org/wiki/Patricia_Schroeder
Patricia Velasquez	http://en.wikipedia.org/wiki/Patricia_Velasquez
Patricia Williams	http://en.wikipedia.org/wiki/Patricia_Williams
Patrick Adiarte	http://en.wikipedia.org/wiki/Patrick_Adiarte
Patrick Dempsey	http://en.wikipedia.org/wiki/Patrick_Dempsey
Patrick Duffy	http://en.wikipedia.org/wiki/Patrick_Duffy
Patrick Ewing	http://en.wikipedia.org/wiki/Patrick_Ewing
Patrick Fugit	http://en.wikipedia.org/wiki/Patrick_Fugit
Patrick Hamilton	http://en.wikipedia.org/wiki/Patrick_Hamilton_(writer)
Patrick Hamilton	http://en.wikipedia.org/wiki/Patrick_Hamilton_(martyr)
Patrick Henry	http://en.wikipedia.org/wiki/Patrick_Henry
Patrick Hillery	http://en.wikipedia.org/wiki/Patrick_Hillery
Patrick J. Fitzgerald	http://en.wikipedia.org/wiki/Patrick_J._Fitzgerald
Patrick J. Hurley	http://en.wikipedia.org/wiki/Patrick_J._Hurley
Patrick J. Moore	http://en.wikipedia.org/wiki/Patrick_J._Moore
Patrick Joseph Kennedy	http://en.wikipedia.org/wiki/Patrick_Joseph_Kennedy
Patrick Kroupa	http://en.wikipedia.org/wiki/Patrick_Kroupa
Patrick Leahy	http://en.wikipedia.org/wiki/Patrick_Leahy
Patrick Leahy	http://en.wikipedia.org/wiki/Patrick_Leahy
Patrick Lichfield	http://en.wikipedia.org/wiki/Patrick_Lichfield
Patrick M. Hughes	http://en.wikipedia.org/wiki/Patrick_M._Hughes
Patrick Macnee	http://en.wikipedia.org/wiki/Patrick_Macnee
Patrick Magee	http://en.wikipedia.org/wiki/Patrick_Magee_(actor)
Patrick Manning	http://en.wikipedia.org/wiki/Patrick_Manning
Patrick Marber	http://en.wikipedia.org/wiki/Patrick_Marber
Patrick McGoohan	http://en.wikipedia.org/wiki/Patrick_McGoohan
Patrick McHenry	http://en.wikipedia.org/wiki/Patrick_McHenry
Patrick McLoughlin	http://en.wikipedia.org/wiki/Patrick_McLoughlin
Patrick Mercer	http://en.wikipedia.org/wiki/Patrick_Mercer
Patrick Moore	http://en.wikipedia.org/wiki/Patrick_Moore
Patrick Muldoon	http://en.wikipedia.org/wiki/Patrick_Muldoon
Patrick Murphy	http://en.wikipedia.org/wiki/Patrick_Murphy_(politician)
Patrick Naughton	http://en.wikipedia.org/wiki/Patrick_Naughton
Patrick Noonan	http://en.wikipedia.org/wiki/Patrick_Noonan
Patrick O'Brian	http://en.wikipedia.org/wiki/Patrick_O%27Brian
Patrick O'Neal	http://en.wikipedia.org/wiki/Patrick_O%27Neal
Patrick Stewart	http://en.wikipedia.org/wiki/Patrick_Stewart
Patrick Stump	http://en.wikipedia.org/wiki/Patrick_Stump
Patrick S�skind	http://en.wikipedia.org/wiki/Patrick_S%FCskind
Patrick Swayze	http://en.wikipedia.org/wiki/Patrick_Swayze
Patrick Troughton	http://en.wikipedia.org/wiki/Patrick_Troughton
Patrick Warburton	http://en.wikipedia.org/wiki/Patrick_Warburton
Patrick Wayne	http://en.wikipedia.org/wiki/Patrick_Wayne
Patrick White	http://en.wikipedia.org/wiki/Patrick_White
Patrick Wilson	http://en.wikipedia.org/wiki/Patrick_Wilson_(actor)
Patrick Wilson	http://en.wikipedia.org/wiki/Patrick_Wilson_(musician)
Patrick Woodroffe	http://en.wikipedia.org/wiki/Patrick_Woodroffe
Patsy Cline	http://en.wikipedia.org/wiki/Patsy_Cline
Patsy Kensit	http://en.wikipedia.org/wiki/Patsy_Kensit
Patsy Ramsey	http://en.wikipedia.org/wiki/Patsy_Ramsey
Patsy Rowlands	http://en.wikipedia.org/wiki/Patsy_Rowlands
Patti Davis	http://en.wikipedia.org/wiki/Patti_Davis
Patti LaBelle	http://en.wikipedia.org/wiki/Patti_LaBelle
Patti LuPone	http://en.wikipedia.org/wiki/Patti_LuPone
Patti Page	http://en.wikipedia.org/wiki/Patti_Page
Patti Smith	http://en.wikipedia.org/wiki/Patti_Smith
Patton Oswalt	http://en.wikipedia.org/wiki/Patton_Oswalt
Patty Andrews	http://en.wikipedia.org/wiki/Patty_Andrews
Patty Duke	http://en.wikipedia.org/wiki/Patty_Duke
Patty Hearst	http://en.wikipedia.org/wiki/Patty_Hearst
Patty Loveless	http://en.wikipedia.org/wiki/Patty_Loveless
Patty Murray	http://en.wikipedia.org/wiki/Patty_Murray
Patty Smyth	http://en.wikipedia.org/wiki/Patty_Smyth
Patty Stonesifer	http://en.wikipedia.org/wiki/Patty_Stonesifer
Paul A. Baran	http://en.wikipedia.org/wiki/Paul_A._Baran
Paul Ableman	http://en.wikipedia.org/wiki/Paul_Ableman
Paul Allaire	http://en.wikipedia.org/wiki/Paul_Allaire
Paul Allen	http://en.wikipedia.org/wiki/Paul_Allen
Paul Ambrose	http://en.wikipedia.org/wiki/Paul_Ambrose
Paul Anka	http://en.wikipedia.org/wiki/Paul_Anka
Paul Atkinson	http://en.wikipedia.org/wiki/Paul_Atkinson_(guitarist)
Paul Auster	http://en.wikipedia.org/wiki/Paul_Auster
Paul B. Henry	http://en.wikipedia.org/wiki/Paul_B._Henry
Paul Bailey	http://en.wikipedia.org/wiki/Paul_Bailey
Paul Banks	http://en.wikipedia.org/wiki/Paul_Banks
Paul Baran	http://en.wikipedia.org/wiki/Paul_Baran
Paul Begala	http://en.wikipedia.org/wiki/Paul_Begala
Paul Benedict	http://en.wikipedia.org/wiki/Paul_Benedict
Paul Ben-Victor	http://en.wikipedia.org/wiki/Paul_Ben-Victor
Paul Beresford	http://en.wikipedia.org/wiki/Paul_Beresford
Paul Berg	http://en.wikipedia.org/wiki/Paul_Berg
Paul Bernardo	http://en.wikipedia.org/wiki/Paul_Bernardo
Paul Bettany	http://en.wikipedia.org/wiki/Paul_Bettany
Paul Biya	http://en.wikipedia.org/wiki/Paul_Biya
Paul Biyogh� Mba	http://en.wikipedia.org/wiki/Paul_Biyogh%E9_Mba
Paul Blomfield	http://en.wikipedia.org/wiki/Paul_Blomfield
Paul Bostaph	http://en.wikipedia.org/wiki/Paul_Bostaph
Paul Bowles	http://en.wikipedia.org/wiki/Paul_Bowles
Paul Broun	http://en.wikipedia.org/wiki/Paul_Broun
Paul Burstow	http://en.wikipedia.org/wiki/Paul_Burstow
Paul Butterfield	http://en.wikipedia.org/wiki/Paul_Butterfield
Paul Carrack	http://en.wikipedia.org/wiki/Paul_Carrack
Paul Castellano	http://en.wikipedia.org/wiki/Paul_Castellano
Paul Cellucci	http://en.wikipedia.org/wiki/Paul_Cellucci
Paul C�zanne	http://en.wikipedia.org/wiki/Paul_C%E9zanne
Paul Claudel	http://en.wikipedia.org/wiki/Paul_Claudel
Paul Coverdell	http://en.wikipedia.org/wiki/Paul_Coverdell
Paul Cronin	http://en.wikipedia.org/wiki/Paul_W._Cronin
Paul Crouch	http://en.wikipedia.org/wiki/Paul_Crouch
Paul D. Boyer	http://en.wikipedia.org/wiki/Paul_D._Boyer
Paul Daniels	http://en.wikipedia.org/wiki/Paul_Daniels
Paul Darrow	http://en.wikipedia.org/wiki/Paul_Darrow
Paul Delaroche	http://en.wikipedia.org/wiki/Paul_Delaroche
Paul Dinello	http://en.wikipedia.org/wiki/Paul_Dinello
Paul Dirac	http://en.wikipedia.org/wiki/Paul_Dirac
Paul Dooley	http://en.wikipedia.org/wiki/Paul_Dooley
Paul Dukas	http://en.wikipedia.org/wiki/Paul_Dukas
Paul E. Kanjorski	http://en.wikipedia.org/wiki/Paul_E._Kanjorski
Paul Eddington	http://en.wikipedia.org/wiki/Paul_Eddington
Paul Ehrlich	http://en.wikipedia.org/wiki/Paul_Ehrlich
Paul Elmer More	http://en.wikipedia.org/wiki/Paul_Elmer_More
Paul �luard	http://en.wikipedia.org/wiki/Paul_%C9luard
Paul Erdos	http://en.wikipedia.org/wiki/Paul_Erdos
Paul F. Tompkins	http://en.wikipedia.org/wiki/Paul_F._Tompkins
Paul Farmer	http://en.wikipedia.org/wiki/Paul_Farmer
Paul Farrelly	http://en.wikipedia.org/wiki/Paul_Farrelly
Paul Flynn	http://en.wikipedia.org/wiki/Paul_Flynn_(politician)
Paul Gascoigne	http://en.wikipedia.org/wiki/Paul_Gascoigne
Paul Gauguin	http://en.wikipedia.org/wiki/Paul_Gauguin
Paul Giamatti	http://en.wikipedia.org/wiki/Paul_Giamatti
Paul Gigot	http://en.wikipedia.org/wiki/Paul_Gigot
Paul Gilbert	http://en.wikipedia.org/wiki/Paul_Gilbert
Paul Gillmor	http://en.wikipedia.org/wiki/Paul_Gillmor
Paul Goggins	http://en.wikipedia.org/wiki/Paul_Goggins
Paul Goodman	http://en.wikipedia.org/wiki/Paul_Goodman_(writer)
Paul Greengrass	http://en.wikipedia.org/wiki/Paul_Greengrass
Paul Gross	http://en.wikipedia.org/wiki/Paul_Gross
Paul Guilfoyle	http://en.wikipedia.org/wiki/Paul_Guilfoyle
Paul H. Allen	http://en.wikipedia.org/wiki/Paul_H._Allen
Paul H. Douglas	http://en.wikipedia.org/wiki/Paul_H._Douglas
Paul Hackett	http://en.wikipedia.org/wiki/Paul_Hackett_(politician)
Paul Hardcastle	http://en.wikipedia.org/wiki/Paul_Hardcastle
Paul Harvey	http://en.wikipedia.org/wiki/Paul_Harvey
Paul Henreid	http://en.wikipedia.org/wiki/Paul_Henreid
Paul Henri d'Estournelles de Constant	http://en.wikipedia.org/wiki/Paul_Henri_d%27Estournelles_de_Constant
Paul Hindemith	http://en.wikipedia.org/wiki/Paul_Hindemith
Paul Hodes	http://en.wikipedia.org/wiki/Paul_Hodes
Paul Hogan	http://en.wikipedia.org/wiki/Paul_Hogan
Paul Horgan	http://en.wikipedia.org/wiki/Paul_Horgan
Paul J. Crutzen	http://en.wikipedia.org/wiki/Paul_J._Crutzen
Paul J. Flory	http://en.wikipedia.org/wiki/Paul_J._Flory
Paul Kagame	http://en.wikipedia.org/wiki/Paul_Kagame
Paul Kammerer	http://en.wikipedia.org/wiki/Paul_Kammerer
Paul Kangas	http://en.wikipedia.org/wiki/Paul_Kangas
Paul Kanjorski	http://en.wikipedia.org/wiki/Paul_Kanjorski
Paul Kantner	http://en.wikipedia.org/wiki/Paul_Kantner
Paul Karrer	http://en.wikipedia.org/wiki/Paul_Karrer
Paul Keating	http://en.wikipedia.org/wiki/Paul_Keating
Paul Klee	http://en.wikipedia.org/wiki/Paul_Klee
Paul Krassner	http://en.wikipedia.org/wiki/Paul_Krassner
Paul Krugman	http://en.wikipedia.org/wiki/Paul_Krugman
Paul Kurtz	http://en.wikipedia.org/wiki/Paul_Kurtz
Paul Langevin	http://en.wikipedia.org/wiki/Paul_Langevin
Paul Laurence Dunbar	http://en.wikipedia.org/wiki/Paul_Laurence_Dunbar
Paul Laxalt	http://en.wikipedia.org/wiki/Paul_Laxalt
Paul Laxalt	http://en.wikipedia.org/wiki/Paul_Laxalt
Paul Le Mat	http://en.wikipedia.org/wiki/Paul_Le_Mat
Paul Lukas	http://en.wikipedia.org/wiki/Paul_Lukas
Paul Lynde	http://en.wikipedia.org/wiki/Paul_Lynde
Paul Lytton	http://en.wikipedia.org/wiki/Paul_Lytton
Paul Maguire	http://en.wikipedia.org/wiki/Paul_Maguire
Paul Martin	http://en.wikipedia.org/wiki/Paul_Martin
Paul Maynard	http://en.wikipedia.org/wiki/Paul_Maynard
Paul Mazursky	http://en.wikipedia.org/wiki/Paul_Mazursky
Paul McCartney	http://en.wikipedia.org/wiki/Paul_McCartney
Paul Meier	http://en.wikipedia.org/wiki/Paul_Meier
Paul Michael Glaser	http://en.wikipedia.org/wiki/Paul_Michael_Glaser
Paul Molitor	http://en.wikipedia.org/wiki/Paul_Molitor
Paul Mooney	http://en.wikipedia.org/wiki/Paul_Mooney_(comedian)
Paul Muldoon	http://en.wikipedia.org/wiki/Paul_Muldoon
Paul Muni	http://en.wikipedia.org/wiki/Paul_Muni
Paul Murphy	http://en.wikipedia.org/wiki/Paul_Murphy_(politician)
Paul Newman	http://en.wikipedia.org/wiki/Paul_Newman
Paul Oakenfold	http://en.wikipedia.org/wiki/Paul_Oakenfold
Paul O'Grady	http://en.wikipedia.org/wiki/Paul_O%27Grady
Paul O'Neill	http://en.wikipedia.org/wiki/Paul_O'Neill_(businessman)
Paul Peter Ewald	http://en.wikipedia.org/wiki/Paul_Peter_Ewald
Paul Petersen	http://en.wikipedia.org/wiki/Paul_Petersen
Paul Pierce	http://en.wikipedia.org/wiki/Paul_Pierce
Paul Prudhomme	http://en.wikipedia.org/wiki/Paul_Prudhomme
Paul R. Ehrlich	http://en.wikipedia.org/wiki/Paul_R._Ehrlich
Paul Reiser	http://en.wikipedia.org/wiki/Paul_Reiser
Paul Reubens	http://en.wikipedia.org/wiki/Paul_Reubens
Paul Revere	http://en.wikipedia.org/wiki/Paul_Revere_&_the_Raiders
Paul Revere	http://en.wikipedia.org/wiki/Paul_Revere
Paul Robeson	http://en.wikipedia.org/wiki/Paul_Robeson
Paul Rodgers	http://en.wikipedia.org/wiki/Paul_Rodgers
Paul Rodriguez	http://en.wikipedia.org/wiki/Paul_Rodriguez
Paul Rudd	http://en.wikipedia.org/wiki/Paul_Rudd
Paul Rudolph	http://en.wikipedia.org/wiki/Paul_Rudolph_(architect)
Paul Ryan	http://en.wikipedia.org/wiki/Paul_Ryan_(politician)
Paul S. Sarbanes	http://en.wikipedia.org/wiki/Paul_S._Sarbanes
Paul S. Trible, Jr.	http://en.wikipedia.org/wiki/Paul_S._Trible%2C_Jr.
Paul Sabatier	http://en.wikipedia.org/wiki/Paul_Sabatier_(chemist)
Paul Samuelson	http://en.wikipedia.org/wiki/Paul_Samuelson
Paul Sarbanes	http://en.wikipedia.org/wiki/Paul_Sarbanes
Paul Schrader	http://en.wikipedia.org/wiki/Paul_Schrader
Paul Scofield	http://en.wikipedia.org/wiki/Paul_Scofield
Paul Scott	http://en.wikipedia.org/wiki/Paul_Mark_Scott
Paul Shaffer	http://en.wikipedia.org/wiki/Paul_Shaffer
Paul Shanley	http://en.wikipedia.org/wiki/Paul_Shanley
Paul Simon	http://en.wikipedia.org/wiki/Paul_Simon
Paul Simon	http://en.wikipedia.org/wiki/Paul_Simon
Paul Sorvino	http://en.wikipedia.org/wiki/Paul_Sorvino
Paul Stanley	http://en.wikipedia.org/wiki/Paul_Stanley
Paul Stookey	http://en.wikipedia.org/wiki/Paul_Stookey
Paul Tagliabue	http://en.wikipedia.org/wiki/Paul_Tagliabue
Paul Theroux	http://en.wikipedia.org/wiki/Paul_Theroux
Paul Thomas	http://en.wikipedia.org/wiki/Paul_Thomas_(bassist)
Paul Thomas Anderson	http://en.wikipedia.org/wiki/Paul_Thomas_Anderson
Paul Tibbets	http://en.wikipedia.org/wiki/Paul_Tibbets
Paul Tillich	http://en.wikipedia.org/wiki/Paul_Tillich
Paul Tonko	http://en.wikipedia.org/wiki/Paul_Tonko
Paul Tsongas	http://en.wikipedia.org/wiki/Paul_Tsongas
Paul Uppal	http://en.wikipedia.org/wiki/Paul_Uppal
Paul Val�ry	http://en.wikipedia.org/wiki/Paul_Val%E9ry
Paul Verhoeven	http://en.wikipedia.org/wiki/Paul_Verhoeven
Paul Verlaine	http://en.wikipedia.org/wiki/Paul_Verlaine
Paul VI	http://en.wikipedia.org/wiki/Paul_VI
Paul Volcker	http://en.wikipedia.org/wiki/Paul_Volcker
Paul von Heyse	http://en.wikipedia.org/wiki/Paul_von_Heyse
Paul von Hindenburg	http://en.wikipedia.org/wiki/Paul_von_Hindenburg
Paul W.S. Anderson	http://en.wikipedia.org/wiki/Paul_W.S._Anderson
Paul Walker	http://en.wikipedia.org/wiki/Paul_Walker
Paul Wall	http://en.wikipedia.org/wiki/Paul_Wall
Paul Watson	http://en.wikipedia.org/wiki/Paul_Watson
Paul Weller	http://en.wikipedia.org/wiki/Paul_Weller
Paul Wellstone	http://en.wikipedia.org/wiki/Paul_Wellstone
Paul Westerberg	http://en.wikipedia.org/wiki/Paul_Westerberg
Paul Westhead	http://en.wikipedia.org/wiki/Paul_Westhead
Paul Weyrich	http://en.wikipedia.org/wiki/Paul_Weyrich
Paul Williams	http://en.wikipedia.org/wiki/Paul_Williams_(songwriter)
Paul Williams	http://en.wikipedia.org/wiki/Paul_Williams_(The_Temptations)
Paul Winchell	http://en.wikipedia.org/wiki/Paul_Winchell
Paul Winfield	http://en.wikipedia.org/wiki/Paul_Winfield
Paul Wolfowitz	http://en.wikipedia.org/wiki/Paul_Wolfowitz
Paul X. Kelley	http://en.wikipedia.org/wiki/Paul_X._Kelley
Paul Young	http://en.wikipedia.org/wiki/Paul_Young
Paul Zindel	http://en.wikipedia.org/wiki/Paul_Zindel
Paula Abdul	http://en.wikipedia.org/wiki/Paula_Abdul
Paula Cole	http://en.wikipedia.org/wiki/Paula_Cole
Paula Hawkins	http://en.wikipedia.org/wiki/Paula_Hawkins
Paula Jones	http://en.wikipedia.org/wiki/Paula_Jones
Paula Marshall	http://en.wikipedia.org/wiki/Paula_Marshall
Paula Poundstone	http://en.wikipedia.org/wiki/Paula_Poundstone
Paula Prentiss	http://en.wikipedia.org/wiki/Paula_Prentiss
Paula Radcliffe	http://en.wikipedia.org/wiki/Paula_Radcliffe
Paula Yates	http://en.wikipedia.org/wiki/Paula_Yates
Paula Zahn	http://en.wikipedia.org/wiki/Paula_Zahn
Paule Marshall	http://en.wikipedia.org/wiki/Paule_Marshall
Paulette Goddard	http://en.wikipedia.org/wiki/Paulette_Goddard
Pauley Perrette	http://en.wikipedia.org/wiki/Pauley_Perrette
Paulina Porizkova	http://en.wikipedia.org/wiki/Paulina_Porizkova
Paulina Rubio	http://en.wikipedia.org/wiki/Paulina_Rubio
Pauline Borghese	http://en.wikipedia.org/wiki/Pauline_Borghese
Pauline Frederick	http://en.wikipedia.org/wiki/Pauline_Frederick
Pauline Frederick	http://en.wikipedia.org/wiki/Pauline_Frederick
Pauline Latham	http://en.wikipedia.org/wiki/Pauline_Latham
Pauline Oliveros	http://en.wikipedia.org/wiki/Pauline_Oliveros
Pauline R�age	http://en.wikipedia.org/wiki/Pauline_R%E9age
Paulo Costanzo	http://en.wikipedia.org/wiki/Paulo_Costanzo
Pauly Shore	http://en.wikipedia.org/wiki/Pauly_Shore
Pavel A. Cherenkov	http://en.wikipedia.org/wiki/Pavel_A._Cherenkov
Pavel Nedved	http://en.wikipedia.org/wiki/Pavel_Nedved
Paz Vega	http://en.wikipedia.org/wiki/Paz_Vega
Peabo Bryson	http://en.wikipedia.org/wiki/Peabo_Bryson
Pearl Bailey	http://en.wikipedia.org/wiki/Pearl_Bailey
Pearl S. Buck	http://en.wikipedia.org/wiki/Pearl_S._Buck
Pearl White	http://en.wikipedia.org/wiki/Pearl_White
Pedro Almod�var	http://en.wikipedia.org/wiki/Pedro_Almod%F3var
Pedro Alonzo Lopez	http://en.wikipedia.org/wiki/Pedro_Alonzo_Lopez
Pedro Bloch	http://en.wikipedia.org/wiki/Pedro_Bloch
Pedro Calder�n de la Barca	http://en.wikipedia.org/wiki/Pedro_Calder%F3n_de_la_Barca
Pedro de Alvarado	http://en.wikipedia.org/wiki/Pedro_de_Alvarado
Pedro II	http://en.wikipedia.org/wiki/Pedro_II_of_Brazil
Pedro Lascurain	http://en.wikipedia.org/wiki/Pedro_Lascurain
Pedro Lazaga	http://en.wikipedia.org/wiki/Pedro_Lazaga
Pedro Martinez	http://en.wikipedia.org/wiki/Pedro_Martinez
Pedro Men�ndez de Avil�s	http://en.wikipedia.org/wiki/Pedro_Men%E9ndez_de_Avil%E9s
Pedro Pablo Kuczynski	http://en.wikipedia.org/wiki/Pedro_Pablo_Kuczynski
Pedro Pires	http://en.wikipedia.org/wiki/Pedro_Pires
Pedro Salinas	http://en.wikipedia.org/wiki/Pedro_Salinas
Pedro Santana Lopes	http://en.wikipedia.org/wiki/Pedro_Santana_Lopes
Pedro the Cruel	http://en.wikipedia.org/wiki/Pedro_the_Cruel
Pee Wee Reese	http://en.wikipedia.org/wiki/Pee_Wee_Reese
Peg Phillips	http://en.wikipedia.org/wiki/Peg_Phillips
Peggy Ashcroft	http://en.wikipedia.org/wiki/Peggy_Ashcroft
Peggy Cass	http://en.wikipedia.org/wiki/Peggy_Cass
Peggy Fleming	http://en.wikipedia.org/wiki/Peggy_Fleming
Peggy Lee	http://en.wikipedia.org/wiki/Peggy_Lee
Peggy Lipton	http://en.wikipedia.org/wiki/Peggy_Lipton
Peggy Mount	http://en.wikipedia.org/wiki/Peggy_Mount
Peggy Noonan	http://en.wikipedia.org/wiki/Peggy_Noonan
Pehr Gyllenhammar	http://en.wikipedia.org/wiki/Pehr_Gyllenhammar
Pele	http://en.wikipedia.org/wiki/Pele
Penelope Ann Miller	http://en.wikipedia.org/wiki/Penelope_Ann_Miller
Penelope Cruz	http://en.wikipedia.org/wiki/Penelope_Cruz
Penelope Fitzgerald	http://en.wikipedia.org/wiki/Penelope_Fitzgerald
Penelope Keith	http://en.wikipedia.org/wiki/Penelope_Keith
Penelope Lively	http://en.wikipedia.org/wiki/Penelope_Lively
Penelope Spheeris	http://en.wikipedia.org/wiki/Penelope_Spheeris
Penn Jillette	http://en.wikipedia.org/wiki/Penn_Jillette
Penny Johnson Jerald	http://en.wikipedia.org/wiki/Penny_Johnson_Jerald
Penny Marshall	http://en.wikipedia.org/wiki/Penny_Marshall
Penny Mordaunt	http://en.wikipedia.org/wiki/Penny_Mordaunt
Per Aage Brandt	http://en.wikipedia.org/wiki/Per_Aage_Brandt
Percival Lowell	http://en.wikipedia.org/wiki/Percival_Lowell
Percy Bysshe Shelley	http://en.wikipedia.org/wiki/Percy_Bysshe_Shelley
Percy Grainger	http://en.wikipedia.org/wiki/Percy_Grainger
Percy MacKaye	http://en.wikipedia.org/wiki/Percy_MacKaye
Percy Sledge	http://en.wikipedia.org/wiki/Percy_Sledge
Percy Williams Bridgman	http://en.wikipedia.org/wiki/Percy_Williams_Bridgman
Perez Prado	http://en.wikipedia.org/wiki/Perez_Prado
Peri Gilpin	http://en.wikipedia.org/wiki/Peri_Gilpin
Perino del Vaga	http://en.wikipedia.org/wiki/Perino_del_Vaga
Perkin Warbeck	http://en.wikipedia.org/wiki/Perkin_Warbeck
Pernell Roberts	http://en.wikipedia.org/wiki/Pernell_Roberts
Pero Bukejlovic	http://en.wikipedia.org/wiki/Pero_Bukejlovic
Perry Christie	http://en.wikipedia.org/wiki/Perry_Christie
Perry Como	http://en.wikipedia.org/wiki/Perry_Como
Perry Farrell	http://en.wikipedia.org/wiki/Perry_Farrell
Perry King	http://en.wikipedia.org/wiki/Perry_King
Perry Miller	http://en.wikipedia.org/wiki/Perry_Miller
Persia White	http://en.wikipedia.org/wiki/Persia_White
Pervez Musharraf	http://en.wikipedia.org/wiki/Pervez_Musharraf
Pervez Musharraf	http://en.wikipedia.org/wiki/Pervez_Musharraf
Peta Wilson	http://en.wikipedia.org/wiki/Peta_Wilson
Pete Best	http://en.wikipedia.org/wiki/Pete_Best
Pete Burns	http://en.wikipedia.org/wiki/Pete_Burns
Pete Conrad	http://en.wikipedia.org/wiki/Pete_Conrad
Pete Coors	http://en.wikipedia.org/wiki/Pete_Coors
Pete Doherty	http://en.wikipedia.org/wiki/Pete_Doherty
Pete Domenici	http://en.wikipedia.org/wiki/Pete_Domenici
Pete du Pont	http://en.wikipedia.org/wiki/Pete_du_Pont
Pete Hamill	http://en.wikipedia.org/wiki/Pete_Hamill
Pete Hoekstra	http://en.wikipedia.org/wiki/Pete_Hoekstra
Pete King	http://en.wikipedia.org/wiki/Peter_T._King
Pete Maravich	http://en.wikipedia.org/wiki/Pete_Maravich
Pete McCloskey	http://en.wikipedia.org/wiki/Pete_McCloskey
Pete Olson	http://en.wikipedia.org/wiki/Pete_Olson
Pete Quaife	http://en.wikipedia.org/wiki/Pete_Quaife
Pete Rose	http://en.wikipedia.org/wiki/Pete_Rose
Pete Rozelle	http://en.wikipedia.org/wiki/Pete_Rozelle
Pete Sampras	http://en.wikipedia.org/wiki/Pete_Sampras
Pete Seeger	http://en.wikipedia.org/wiki/Pete_Seeger
Pete Sessions	http://en.wikipedia.org/wiki/Pete_Sessions
Pete Shelley	http://en.wikipedia.org/wiki/Pete_Shelley
Pete Stark	http://en.wikipedia.org/wiki/Pete_Stark
Pete Stark	http://en.wikipedia.org/wiki/Pete_Stark
Pete Townshend	http://en.wikipedia.org/wiki/Pete_Townshend
Pete V. Domenici	http://en.wikipedia.org/wiki/Pete_V._Domenici
Pete Wiggs	http://en.wikipedia.org/wiki/Pete_Wiggs
Pete Williams	http://en.wikipedia.org/wiki/Harrison_A._Williams
Pete Wilson	http://en.wikipedia.org/wiki/Pete_Wilson
Pete Wilson	http://en.wikipedia.org/wiki/Pete_Wilson
Pete Wilson	http://en.wikipedia.org/wiki/Pete_Wilson_(broadcaster)
Pete Wishart	http://en.wikipedia.org/wiki/Pete_Wishart
Peter Abbay	http://en.wikipedia.org/wiki/Peter_Abbay
Peter Abelard	http://en.wikipedia.org/wiki/Peter_Abelard
Peter Abrahams	http://en.wikipedia.org/wiki/Peter_Abrahams
Peter Ackroyd	http://en.wikipedia.org/wiki/Peter_Ackroyd
Peter Agre	http://en.wikipedia.org/wiki/Peter_Agre
Peter Akinola	http://en.wikipedia.org/wiki/Peter_Akinola
Peter Aldous	http://en.wikipedia.org/wiki/Peter_Aldous
Peter Allen	http://en.wikipedia.org/wiki/Peter_Allen_(composer)
Peter Allen	http://en.wikipedia.org/wiki/Peter_Allen
Peter Andr�	http://en.wikipedia.org/wiki/Peter_Andr%E9
Peter Andreas Hansen	http://en.wikipedia.org/wiki/Peter_Andreas_Hansen
Peter Arnett	http://en.wikipedia.org/wiki/Peter_Arnett
Peter Asher	http://en.wikipedia.org/wiki/Peter_Asher
Peter Bagge	http://en.wikipedia.org/wiki/Peter_Bagge
Peter Banks	http://en.wikipedia.org/wiki/Peter_Banks
Peter Bart	http://en.wikipedia.org/wiki/Peter_Bart
Peter Behrens	http://en.wikipedia.org/wiki/Peter_Behrens
Peter Benchley	http://en.wikipedia.org/wiki/Peter_Benchley
Peter Benenson	http://en.wikipedia.org/wiki/Peter_Benenson
Peter Berg	http://en.wikipedia.org/wiki/Peter_Berg
Peter Billingsley	http://en.wikipedia.org/wiki/Peter_Billingsley
Peter Black	http://en.wikipedia.org/wiki/Peter_Black_(Australian_politician)
Peter Blegvad	http://en.wikipedia.org/wiki/Peter_Blegvad
Peter Bogdanovich	http://en.wikipedia.org/wiki/Peter_Bogdanovich
Peter Bone	http://en.wikipedia.org/wiki/Peter_Bone
Peter Bonerz	http://en.wikipedia.org/wiki/Peter_Bonerz
Peter Bottomley	http://en.wikipedia.org/wiki/Peter_Bottomley
Peter Boyle	http://en.wikipedia.org/wiki/Peter_Boyle
Peter Breck	http://en.wikipedia.org/wiki/Peter_Breck
Peter Brock	http://en.wikipedia.org/wiki/Peter_Brock
Peter Brook	http://en.wikipedia.org/wiki/Peter_Brook
Peter Buck	http://en.wikipedia.org/wiki/Peter_Buck
Peter Burwash	http://en.wikipedia.org/wiki/Peter_Burwash
Peter Camejo	http://en.wikipedia.org/wiki/Peter_Camejo
Peter Caruana	http://en.wikipedia.org/wiki/Peter_Caruana
Peter Cetera	http://en.wikipedia.org/wiki/Peter_Cetera
Peter Christopherson	http://en.wikipedia.org/wiki/Peter_Christopherson
Peter Cook	http://en.wikipedia.org/wiki/Peter_Cook
Peter Coyote	http://en.wikipedia.org/wiki/Peter_Coyote
Peter Criss	http://en.wikipedia.org/wiki/Peter_Criss
Peter Cushing	http://en.wikipedia.org/wiki/Peter_Cushing
Peter D. Ouspensky	http://en.wikipedia.org/wiki/Peter_D._Ouspensky
Peter Davison	http://en.wikipedia.org/wiki/Peter_Davison
Peter Debye	http://en.wikipedia.org/wiki/Peter_Debye
Peter DeFazio	http://en.wikipedia.org/wiki/Peter_DeFazio
Peter DeLuise	http://en.wikipedia.org/wiki/Peter_DeLuise
Peter Deutsch	http://en.wikipedia.org/wiki/Peter_Deutsch
Peter Diamandis	http://en.wikipedia.org/wiki/Peter_Diamandis
Peter Dinklage	http://en.wikipedia.org/wiki/Peter_Dinklage
Peter Drucker	http://en.wikipedia.org/wiki/Peter_Drucker
Peter Facinelli	http://en.wikipedia.org/wiki/Peter_Facinelli
Peter Falk	http://en.wikipedia.org/wiki/Peter_Falk
Peter Farrelly	http://en.wikipedia.org/wiki/Peter_Farrelly
Peter Finch	http://en.wikipedia.org/wiki/Peter_Finch
Peter Fitzgerald	http://en.wikipedia.org/wiki/Peter_Fitzgerald_(politician)
Peter Fonda	http://en.wikipedia.org/wiki/Peter_Fonda
Peter Frampton	http://en.wikipedia.org/wiki/Peter_Frampton
Peter Frelinghuysen, Jr.	http://en.wikipedia.org/wiki/Peter_Frelinghuysen%2C_Jr.
Peter G. Peterson	http://en.wikipedia.org/wiki/Peter_G._Peterson
Peter Gabriel	http://en.wikipedia.org/wiki/Peter_Gabriel
Peter Galbraith	http://en.wikipedia.org/wiki/Peter_Galbraith
Peter Gallagher	http://en.wikipedia.org/wiki/Peter_Gallagher
Peter Garrett	http://en.wikipedia.org/wiki/Peter_Garrett
Peter Gay	http://en.wikipedia.org/wiki/Peter_Gay
Peter Giles	http://en.wikipedia.org/wiki/Peter_Giles_(musician)
Peter Gotti	http://en.wikipedia.org/wiki/Peter_Gotti
Peter Graves	http://en.wikipedia.org/wiki/Peter_Graves_(actor)
Peter Green	http://en.wikipedia.org/wiki/Peter_Green_(musician)
Peter Greenaway	http://en.wikipedia.org/wiki/Peter_Greenaway
Peter Guthrie Tait	http://en.wikipedia.org/wiki/Peter_Guthrie_Tait
Peter H. Kostmayer	http://en.wikipedia.org/wiki/Peter_H._Kostmayer
Peter Hain	http://en.wikipedia.org/wiki/Peter_Hain
Peter Hall	http://en.wikipedia.org/wiki/Peter_W._Hall
Peter Hermann	http://en.wikipedia.org/wiki/Peter_Hermann
Peter Hewitt	http://en.wikipedia.org/wiki/Peter_Hewitt_(film_director)
Peter Hook	http://en.wikipedia.org/wiki/Peter_Hook
Peter Horton	http://en.wikipedia.org/wiki/Peter_Horton
Peter Hyams	http://en.wikipedia.org/wiki/Peter_Hyams
Peter Ilyich Tchaikovsky	http://en.wikipedia.org/wiki/Peter_Ilyich_Tchaikovsky
Peter J. Brennan	http://en.wikipedia.org/wiki/Peter_J._Brennan
Peter J. Visclosky	http://en.wikipedia.org/wiki/Peter_J._Visclosky
Peter Jackson	http://en.wikipedia.org/wiki/Peter_Jackson
Peter Jennings	http://en.wikipedia.org/wiki/Peter_Jennings
Peter Jurasik	http://en.wikipedia.org/wiki/Peter_Jurasik
Peter Krause	http://en.wikipedia.org/wiki/Peter_Krause
Peter Kropotkin	http://en.wikipedia.org/wiki/Peter_Kropotkin
Peter Kruder	http://en.wikipedia.org/wiki/Peter_Kruder
Peter Lawford	http://en.wikipedia.org/wiki/Peter_Lawford
Peter Lilley	http://en.wikipedia.org/wiki/Peter_Lilley
Peter Lombard	http://en.wikipedia.org/wiki/Peter_Lombard
Peter Lorre	http://en.wikipedia.org/wiki/Peter_Lorre
Peter Luff	http://en.wikipedia.org/wiki/Peter_Luff
Peter Maas	http://en.wikipedia.org/wiki/Peter_Maas
Peter Mark Roget	http://en.wikipedia.org/wiki/Peter_Mark_Roget
Peter Marshall	http://en.wikipedia.org/wiki/Peter_Marshall_(U.S._entertainer)
Peter Matthiessen	http://en.wikipedia.org/wiki/Peter_Matthiessen
Peter Max	http://en.wikipedia.org/wiki/Peter_Max
Peter Mayhew	http://en.wikipedia.org/wiki/Peter_Mayhew
Peter Medawar	http://en.wikipedia.org/wiki/Peter_Medawar
Peter Mitchell	http://en.wikipedia.org/wiki/Peter_D._Mitchell
Peter Munk	http://en.wikipedia.org/wiki/Peter_Munk
Peter Murphy	http://en.wikipedia.org/wiki/Peter_Murphy_(musician)
Peter Noone	http://en.wikipedia.org/wiki/Peter_Noone
Peter Norton	http://en.wikipedia.org/wiki/Peter_Norton
Peter of Savoy	http://en.wikipedia.org/wiki/Peter_II_of_Savoy
Peter Oliver	http://en.wikipedia.org/wiki/Peter_Oliver_(painter)
Peter Orlovsky	http://en.wikipedia.org/wiki/Peter_Orlovsky
Peter O'Toole	http://en.wikipedia.org/wiki/Peter_O%27Toole
Peter Pace	http://en.wikipedia.org/wiki/Peter_Pace
Peter Paige	http://en.wikipedia.org/wiki/Peter_Paige
Peter Paul Rubens	http://en.wikipedia.org/wiki/Peter_Paul_Rubens
Peter Popoff	http://en.wikipedia.org/wiki/Peter_Popoff
Peter Riegert	http://en.wikipedia.org/wiki/Peter_Riegert
Peter Roskam	http://en.wikipedia.org/wiki/Peter_Roskam
Peter Sarsgaard	http://en.wikipedia.org/wiki/Peter_Sarsgaard
Peter Schmeichel	http://en.wikipedia.org/wiki/Peter_Schmeichel
Peter Scolari	http://en.wikipedia.org/wiki/Peter_Scolari
Peter Segal	http://en.wikipedia.org/wiki/Peter_Segal
Peter Sellers	http://en.wikipedia.org/wiki/Peter_Sellers
Peter Shaffer	http://en.wikipedia.org/wiki/Peter_Shaffer
Peter Singer	http://en.wikipedia.org/wiki/Peter_Singer
Peter Sotos	http://en.wikipedia.org/wiki/Peter_Sotos
Peter Soulsby	http://en.wikipedia.org/wiki/Peter_Soulsby
Peter Steele	http://en.wikipedia.org/wiki/Peter_Steele
Peter Stormare	http://en.wikipedia.org/wiki/Peter_Stormare
Peter Straub	http://en.wikipedia.org/wiki/Peter_Straub
Peter Strauss	http://en.wikipedia.org/wiki/Peter_Strauss
Peter Struck	http://en.wikipedia.org/wiki/Peter_Struck
Peter Stuyvesant	http://en.wikipedia.org/wiki/Peter_Stuyvesant
Peter Sutcliffe	http://en.wikipedia.org/wiki/Peter_Sutcliffe
Peter Sutherland	http://en.wikipedia.org/wiki/Peter_Sutherland
Peter Tapsell	http://en.wikipedia.org/wiki/Peter_Tapsell_(UK_politician)
Peter Taylor	http://en.wikipedia.org/wiki/Peter_Matthew_Hillsman_Taylor
Peter the Great	http://en.wikipedia.org/wiki/Peter_the_Great
Peter the Hermit	http://en.wikipedia.org/wiki/Peter_the_Hermit
Peter Thomson	http://en.wikipedia.org/wiki/Peter_Thomson_(Australian_golfer)
Peter Tomarken	http://en.wikipedia.org/wiki/Peter_Tomarken
Peter Tork	http://en.wikipedia.org/wiki/Peter_Tork
Peter Tosh	http://en.wikipedia.org/wiki/Peter_Tosh
Peter Ueberroth	http://en.wikipedia.org/wiki/Peter_Ueberroth
Peter Ustinov	http://en.wikipedia.org/wiki/Peter_Ustinov
Peter Viereck	http://en.wikipedia.org/wiki/Peter_Viereck
Peter Visclosky	http://en.wikipedia.org/wiki/Peter_Visclosky
Peter W. Rodino, Jr.	http://en.wikipedia.org/wiki/Peter_W._Rodino%2C_Jr.
Peter Weir	http://en.wikipedia.org/wiki/Peter_Weir
Peter Welch	http://en.wikipedia.org/wiki/Peter_Welch
Peter Weller	http://en.wikipedia.org/wiki/Peter_Weller
Peter Wentz	http://en.wikipedia.org/wiki/Peter_Wentz
Peter Yarrow	http://en.wikipedia.org/wiki/Peter_Yarrow
Peter Yates	http://en.wikipedia.org/wiki/Peter_Yates
Petey Pablo	http://en.wikipedia.org/wiki/Petey_Pablo
Petra Haden	http://en.wikipedia.org/wiki/Petra_Haden
Petroleum V. Nasby	http://en.wikipedia.org/wiki/Petroleum_V._Nasby
Petronius Arbiter	http://en.wikipedia.org/wiki/Petronius_Arbiter
Petula Clark	http://en.wikipedia.org/wiki/Petula_Clark
Peyton Manning	http://en.wikipedia.org/wiki/Peyton_Manning
Peyton Randolph	http://en.wikipedia.org/wiki/Peyton_Randolph
Phan Van Khai	http://en.wikipedia.org/wiki/Phan_Van_Khai
Pharrell Williams	http://en.wikipedia.org/wiki/Pharrell_Williams
Phil Angelides	http://en.wikipedia.org/wiki/Phil_Angelides
Phil Anselmo	http://en.wikipedia.org/wiki/Phil_Anselmo
Phil Bredesen	http://en.wikipedia.org/wiki/Phil_Bredesen
Phil Bredesen	http://en.wikipedia.org/wiki/Phil_Bredesen
Phil Brown	http://en.wikipedia.org/wiki/Phil_Brown_(actor)
Phil Collen	http://en.wikipedia.org/wiki/Phil_Collen
Phil Collins	http://en.wikipedia.org/wiki/Phil_Collins
Phil Crane	http://en.wikipedia.org/wiki/Phil_Crane
Phil Donahue	http://en.wikipedia.org/wiki/Phil_Donahue
Phil English	http://en.wikipedia.org/wiki/Phil_English
Phil Esposito	http://en.wikipedia.org/wiki/Phil_Esposito
Phil Everly	http://en.wikipedia.org/wiki/Phil_Everly
Phil Foglio	http://en.wikipedia.org/wiki/Phil_Foglio
Phil Gingrey	http://en.wikipedia.org/wiki/Phil_Gingrey
Phil Gramm	http://en.wikipedia.org/wiki/Phil_Gramm
Phil Gramm	http://en.wikipedia.org/wiki/Phil_Gramm
Phil Hare	http://en.wikipedia.org/wiki/Phil_Hare
Phil Harris	http://en.wikipedia.org/wiki/Phil_Harris
Phil Hartman	http://en.wikipedia.org/wiki/Phil_Hartman
Phil Hay	http://en.wikipedia.org/wiki/Phil_Hay
Phil Katz	http://en.wikipedia.org/wiki/Phil_Katz
Phil Knight	http://en.wikipedia.org/wiki/Phil_Knight
Phil LaMarr	http://en.wikipedia.org/wiki/Phil_LaMarr
Phil Lesh	http://en.wikipedia.org/wiki/Phil_Lesh
Phil Lynott	http://en.wikipedia.org/wiki/Phil_Lynott
Phil Margera	http://en.wikipedia.org/wiki/Phil_Margera
Phil Mickelson	http://en.wikipedia.org/wiki/Phil_Mickelson
Phil Miller	http://en.wikipedia.org/wiki/Phil_Miller
Phil Ochs	http://en.wikipedia.org/wiki/Phil_Ochs
Phil Rizzuto	http://en.wikipedia.org/wiki/Phil_Rizzuto
Phil Roe	http://en.wikipedia.org/wiki/Phil_Roe
Phil Rudd	http://en.wikipedia.org/wiki/Phil_Rudd
Phil Selway	http://en.wikipedia.org/wiki/Phil_Selway
Phil Silvers	http://en.wikipedia.org/wiki/Phil_Silvers
Phil Spector	http://en.wikipedia.org/wiki/Phil_Spector
Phil Wilson	http://en.wikipedia.org/wiki/Phil_Wilson_(British_politician)
Phil Woolas	http://en.wikipedia.org/wiki/Phil_Woolas
Phil Zimmermann	http://en.wikipedia.org/wiki/Phil_Zimmermann
Philander Knox	http://en.wikipedia.org/wiki/Philander_Knox
Phil�mon Yang	http://en.wikipedia.org/wiki/Phil%E9mon_Yang
Philetas of Cos	http://en.wikipedia.org/wiki/Philetas_of_Cos
Philip Anschutz	http://en.wikipedia.org/wiki/Philip_Anschutz
Philip Bailey	http://en.wikipedia.org/wiki/Philip_Bailey
Philip Bailhache	http://en.wikipedia.org/wiki/Philip_Bailhache
Philip Baker Hall	http://en.wikipedia.org/wiki/Philip_Baker_Hall
Philip Caputo	http://en.wikipedia.org/wiki/Philip_Caputo
Philip Crosby	http://en.wikipedia.org/wiki/Phillip_Crosby
Philip Davies	http://en.wikipedia.org/wiki/Philip_Davies
Philip Dunne	http://en.wikipedia.org/wiki/Philip_Dunne_(politician)
Philip Glass	http://en.wikipedia.org/wiki/Philip_Glass
Philip Greenspun	http://en.wikipedia.org/wiki/Philip_Greenspun
Philip Hammond	http://en.wikipedia.org/wiki/Philip_Hammond
Philip Henry Sheridan	http://en.wikipedia.org/wiki/Philip_Henry_Sheridan
Philip Henslowe	http://en.wikipedia.org/wiki/Philip_Henslowe
Philip Hollobone	http://en.wikipedia.org/wiki/Philip_Hollobone
Philip I	http://en.wikipedia.org/wiki/Philip_I_of_Castile
Philip II	http://en.wikipedia.org/wiki/Philip_II_of_Spain
Philip III	http://en.wikipedia.org/wiki/Philip_III_of_Spain
Philip IV	http://en.wikipedia.org/wiki/Philip_IV_of_Spain
Philip J. Kaplan	http://en.wikipedia.org/wiki/Philip_J._Kaplan
Philip J. Purcell	http://en.wikipedia.org/wiki/Philip_J._Purcell
Philip Jeck	http://en.wikipedia.org/wiki/Philip_Jeck
Philip Johnson	http://en.wikipedia.org/wiki/Philip_Johnson
Philip Jos� Farmer	http://en.wikipedia.org/wiki/Philip_Jos%E9_Farmer
Philip K. Dick	http://en.wikipedia.org/wiki/Philip_K._Dick
Philip Kearny	http://en.wikipedia.org/wiki/Philip_Kearny
Philip Larkin	http://en.wikipedia.org/wiki/Philip_Larkin
Philip Lee	http://en.wikipedia.org/wiki/Phillip_Lee_(politician)
Philip Levine	http://en.wikipedia.org/wiki/Philip_Levine_(poet)
Philip M. Crane	http://en.wikipedia.org/wiki/Philip_M._Crane
Philip M. Klutznick	http://en.wikipedia.org/wiki/Philip_M._Klutznick
Philip Massinger	http://en.wikipedia.org/wiki/Philip_Massinger
Philip McKeon	http://en.wikipedia.org/wiki/Philip_McKeon
Philip Michael Thomas	http://en.wikipedia.org/wiki/Philip_Michael_Thomas
Philip Neri	http://en.wikipedia.org/wiki/Philip_Neri
Philip Noel-Baker	http://en.wikipedia.org/wiki/Philip_Noel-Baker
Philip R. Sharp	http://en.wikipedia.org/wiki/Philip_R._Sharp
Philip Rahv	http://en.wikipedia.org/wiki/Philip_Rahv
Philip Roth	http://en.wikipedia.org/wiki/Philip_Roth
Philip Schuyler	http://en.wikipedia.org/wiki/Philip_Schuyler
Philip Seymour Hoffman	http://en.wikipedia.org/wiki/Philip_Seymour_Hoffman
Philip Stephens	http://en.wikipedia.org/wiki/Philip_Stephens_(journalist)
Philip the Arab	http://en.wikipedia.org/wiki/Philip_the_Arab
Philip V	http://en.wikipedia.org/wiki/Philip_V_of_Spain
Philip W. Anderson	http://en.wikipedia.org/wiki/Philip_W._Anderson
Philip Whalen	http://en.wikipedia.org/wiki/Philip_Whalen
Philip Zelikow	http://en.wikipedia.org/wiki/Philip_Zelikow
Philip Zimbardo	http://en.wikipedia.org/wiki/Philip_Zimbardo
Philipp Lenard	http://en.wikipedia.org/wiki/Philipp_Lenard
Philipp Melanchthon	http://en.wikipedia.org/wiki/Philipp_Melanchthon
Philipp Scheidemann	http://en.wikipedia.org/wiki/Philipp_Scheidemann
Philippa of Hainaut	http://en.wikipedia.org/wiki/Philippa_of_Hainaut
Philippe Busquin	http://en.wikipedia.org/wiki/Philippe_Busquin
Philippe de Champaigne	http://en.wikipedia.org/wiki/Philippe_de_Champaigne
Philippe I	http://en.wikipedia.org/wiki/Philip_I_of_France
Philippe II	http://en.wikipedia.org/wiki/Philip_II_of_France
Philippe II, duc d'Orl�ans	http://en.wikipedia.org/wiki/Philippe_II%2C_duc_d%27Orl%E9ans
Philippe III	http://en.wikipedia.org/wiki/Philippe_III
Philippe IV	http://en.wikipedia.org/wiki/Philippe_IV
Philippe Leroy	http://en.wikipedia.org/wiki/Philippe_Leroy_(actor)
Philippe Noiret	http://en.wikipedia.org/wiki/Philippe_Noiret
Philippe P�tain	http://en.wikipedia.org/wiki/Philippe_P%E9tain
Philippe V	http://en.wikipedia.org/wiki/Philip_V_of_France
Philippe VI	http://en.wikipedia.org/wiki/Philippe_VI
Phill Kline	http://en.wikipedia.org/wiki/Phill_Kline
Phillip Alford	http://en.wikipedia.org/wiki/Phillip_Alford
Phillip Burton	http://en.wikipedia.org/wiki/Phillip_Burton
Phillip Johnson	http://en.wikipedia.org/wiki/Phillip_E._Johnson
Phillip Noyce	http://en.wikipedia.org/wiki/Phillip_Noyce
Phillis Wheatley	http://en.wikipedia.org/wiki/Phillis_Wheatley
Philo Farnsworth	http://en.wikipedia.org/wiki/Philo_Farnsworth
Phoebe Cates	http://en.wikipedia.org/wiki/Phoebe_Cates
Phoebe Snow	http://en.wikipedia.org/wiki/Phoebe_Snow
Phoenix Farrell	http://en.wikipedia.org/wiki/Phoenix_Farrell
Phylicia Rashad	http://en.wikipedia.org/wiki/Phylicia_Rashad
Phylicia Rashad	http://en.wikipedia.org/wiki/Phylicia_Rashad
Phyllis Diller	http://en.wikipedia.org/wiki/Phyllis_Diller
Phyllis Fraser	http://en.wikipedia.org/wiki/Phyllis_Fraser
Phyllis George	http://en.wikipedia.org/wiki/Phyllis_George
Phyllis Hyman	http://en.wikipedia.org/wiki/Phyllis_Hyman
Phyllis McGinley	http://en.wikipedia.org/wiki/Phyllis_McGinley
Phyllis Schlafly	http://en.wikipedia.org/wiki/Phyllis_Schlafly
Pia Zadora	http://en.wikipedia.org/wiki/Pia_Zadora
Pier Angeli	http://en.wikipedia.org/wiki/Pier_Angeli
Pier Luigi Nervi	http://en.wikipedia.org/wiki/Pier_Luigi_Nervi
Pier Paolo Pasolini	http://en.wikipedia.org/wiki/Pier_Paolo_Pasolini
Pierce Brosnan	http://en.wikipedia.org/wiki/Pierce_Brosnan
Piero della Francesca	http://en.wikipedia.org/wiki/Piero_della_Francesca
Piero Umiliani	http://en.wikipedia.org/wiki/Piero_Umiliani
Pierre Akendengue	http://en.wikipedia.org/wiki/Pierre_Akendengue
Pierre Beaumarchais	http://en.wikipedia.org/wiki/Pierre_Beaumarchais
Pierre Belon	http://en.wikipedia.org/wiki/Pierre_Belon
Pierre B�r�govoy	http://en.wikipedia.org/wiki/Pierre_B%E9r%E9govoy
Pierre Berton	http://en.wikipedia.org/wiki/Pierre_Berton
Pierre Bonnard	http://en.wikipedia.org/wiki/Pierre_Bonnard
Pierre Bouguer	http://en.wikipedia.org/wiki/Pierre_Bouguer
Pierre Boulez	http://en.wikipedia.org/wiki/Pierre_Boulez
Pierre Bouvier	http://en.wikipedia.org/wiki/Pierre_Bouvier
Pierre Cardin	http://en.wikipedia.org/wiki/Pierre_Cardin
Pierre Charles L'Enfant	http://en.wikipedia.org/wiki/Pierre_Charles_L%27Enfant
Pierre Charron	http://en.wikipedia.org/wiki/Pierre_Charron
Pierre Choderlos de Laclos	http://en.wikipedia.org/wiki/Pierre_Choderlos_de_Laclos
Pierre Corneille	http://en.wikipedia.org/wiki/Pierre_Corneille
Pierre Curie	http://en.wikipedia.org/wiki/Pierre_Curie
Pierre de Brant�me	http://en.wikipedia.org/wiki/Pierre_de_Brant%F4me
Pierre de Fermat	http://en.wikipedia.org/wiki/Pierre_de_Fermat
Pierre de Ronsard	http://en.wikipedia.org/wiki/Pierre_de_Ronsard
Pierre Dupuy	http://en.wikipedia.org/wiki/Pierre_Dupuy_(scholar)
Pierre Gemayel	http://en.wikipedia.org/wiki/Pierre_Gemayel
Pierre Gustave Toutant Beauregard	http://en.wikipedia.org/wiki/Pierre_Gustave_Toutant_Beauregard
Pierre Henry	http://en.wikipedia.org/wiki/Pierre_Henry
Pierre Janet	http://en.wikipedia.org/wiki/Pierre_Janet
Pierre Janssen	http://en.wikipedia.org/wiki/Pierre_Janssen
Pierre Laval	http://en.wikipedia.org/wiki/Pierre_Laval
Pierre Marivaux	http://en.wikipedia.org/wiki/Pierre_Marivaux
Pierre Nkurunziza	http://en.wikipedia.org/wiki/Pierre_Nkurunziza
Pierre Omidyar	http://en.wikipedia.org/wiki/Pierre_Omidyar
Pierre Pettigrew	http://en.wikipedia.org/wiki/Pierre_Pettigrew
Pierre Poujade	http://en.wikipedia.org/wiki/Pierre_Poujade
Pierre Salinger	http://en.wikipedia.org/wiki/Pierre_Salinger
Pierre Schaeffer	http://en.wikipedia.org/wiki/Pierre_Schaeffer
Pierre Teilhard de Chardin	http://en.wikipedia.org/wiki/Pierre_Teilhard_de_Chardin
Pierre Trudeau	http://en.wikipedia.org/wiki/Pierre_Trudeau
Pierre-Daniel Huet	http://en.wikipedia.org/wiki/Pierre-Daniel_Huet
Pierre-Fran�ois-Xavier de Charlevoix	http://en.wikipedia.org/wiki/Pierre-Fran%E7ois-Xavier_de_Charlevoix
Pierre-Gilles de Gennes	http://en.wikipedia.org/wiki/Pierre-Gilles_de_Gennes
Pierre-Jean David d'Angers	http://en.wikipedia.org/wiki/Pierre-Jean_David_d%27Angers
Pierre-Joseph Desault	http://en.wikipedia.org/wiki/Pierre-Joseph_Desault
Pierre-Louis Moreau de Maupertuis	http://en.wikipedia.org/wiki/Pierre-Louis_Moreau_de_Maupertuis
Pierre-Simon Laplace	http://en.wikipedia.org/wiki/Pierre-Simon_Laplace
Piers Anthony	http://en.wikipedia.org/wiki/Piers_Anthony
Piet Joubert	http://en.wikipedia.org/wiki/Piet_Joubert
Piet Mondrian	http://en.wikipedia.org/wiki/Piet_Mondrian
Pieter Brueghel	http://en.wikipedia.org/wiki/Pieter_Brueghel_the_Elder
Pieter Corneliszoon Hooft	http://en.wikipedia.org/wiki/Pieter_Corneliszoon_Hooft
Pieter de Hooch	http://en.wikipedia.org/wiki/Pieter_de_Hooch
Pieter Zeeman	http://en.wikipedia.org/wiki/Pieter_Zeeman
Pietro Aretino	http://en.wikipedia.org/wiki/Pietro_Aretino
Pietro Cavallini	http://en.wikipedia.org/wiki/Pietro_Cavallini
Pietro Damiani	http://en.wikipedia.org/wiki/Pietro_Damiani
Pietro Longhi	http://en.wikipedia.org/wiki/Pietro_Longhi
Pietro Mascagni	http://en.wikipedia.org/wiki/Pietro_Mascagni
Pim Fortuyn	http://en.wikipedia.org/wiki/Pim_Fortuyn
Pio Tuia	http://en.wikipedia.org/wiki/Pio_Tuia
Pip Pyle	http://en.wikipedia.org/wiki/Pip_Pyle
Piper Laurie	http://en.wikipedia.org/wiki/Piper_Laurie
Piper Perabo	http://en.wikipedia.org/wiki/Piper_Perabo
Pitts Sanborn	http://en.wikipedia.org/wiki/Pitts_Sanborn
Pius VIII	http://en.wikipedia.org/wiki/Pius_VIII
Pius XI	http://en.wikipedia.org/wiki/Pius_XI
Pius XII	http://en.wikipedia.org/wiki/Pius_XII
Placido Domingo	http://en.wikipedia.org/wiki/Placido_Domingo
Pol Pot	http://en.wikipedia.org/wiki/Pol_Pot
Pola Negri	http://en.wikipedia.org/wiki/Pola_Negri
Polidoro Caldara da Caravaggio	http://en.wikipedia.org/wiki/Polidoro_Caldara_da_Caravaggio
Polly Bergen	http://en.wikipedia.org/wiki/Polly_Bergen
Polly Holliday	http://en.wikipedia.org/wiki/Polly_Holliday
Polly Klaas	http://en.wikipedia.org/wiki/Polly_Klaas
Polykarp Kusch	http://en.wikipedia.org/wiki/Polykarp_Kusch
Pope Adrian I	http://en.wikipedia.org/wiki/Pope_Adrian_I
Pope Adrian II	http://en.wikipedia.org/wiki/Pope_Adrian_II
Pope Adrian IV	http://en.wikipedia.org/wiki/Pope_Adrian_IV
Pope Adrian VI	http://en.wikipedia.org/wiki/Pope_Adrian_VI
Pope Agatho	http://en.wikipedia.org/wiki/Pope_Agatho
Pope Alexander II	http://en.wikipedia.org/wiki/Pope_Alexander_II
Pope Alexander III	http://en.wikipedia.org/wiki/Pope_Alexander_III
Pope Alexander V	http://en.wikipedia.org/wiki/Pope_Alexander_V
Pope Alexander VI	http://en.wikipedia.org/wiki/Pope_Alexander_VI
Pope Alexander VII	http://en.wikipedia.org/wiki/Pope_Alexander_VII
Pope Alexander VIII	http://en.wikipedia.org/wiki/Pope_Alexander_VIII
Pope Benedict IX	http://en.wikipedia.org/wiki/Pope_Benedict_IX
Pope Benedict XI	http://en.wikipedia.org/wiki/Pope_Benedict_XI
Pope Benedict XII	http://en.wikipedia.org/wiki/Pope_Benedict_XII
Pope Benedict XIII	http://en.wikipedia.org/wiki/Pope_Benedict_XIII
Pope Benedict XIV	http://en.wikipedia.org/wiki/Pope_Benedict_XIV
Pope Benedict XV	http://en.wikipedia.org/wiki/Pope_Benedict_XV
Pope Benedict XVI	http://en.wikipedia.org/wiki/Pope_Benedict_XVI
Pope Callistus III	http://en.wikipedia.org/wiki/Pope_Callistus_III
Pope Celestine I	http://en.wikipedia.org/wiki/Pope_Celestine_I
Pope Celestine II	http://en.wikipedia.org/wiki/Pope_Celestine_II
Pope Celestine III	http://en.wikipedia.org/wiki/Pope_Celestine_III
Pope Celestine IV	http://en.wikipedia.org/wiki/Pope_Celestine_IV
Pope Celestine V	http://en.wikipedia.org/wiki/Pope_Celestine_V
Pope Clement II	http://en.wikipedia.org/wiki/Pope_Clement_II
Pope Clement III	http://en.wikipedia.org/wiki/Pope_Clement_III
Pope Clement IV	http://en.wikipedia.org/wiki/Pope_Clement_IV
Pope Clement IX	http://en.wikipedia.org/wiki/Pope_Clement_IX
Pope Clement V	http://en.wikipedia.org/wiki/Pope_Clement_V
Pope Clement VI	http://en.wikipedia.org/wiki/Pope_Clement_VI
Pope Clement VII	http://en.wikipedia.org/wiki/Pope_Clement_VII
Pope Clement VIII	http://en.wikipedia.org/wiki/Pope_Clement_VIII
Pope Clement X	http://en.wikipedia.org/wiki/Pope_Clement_X
Pope Clement XI	http://en.wikipedia.org/wiki/Pope_Clement_XI
Pope Clement XII	http://en.wikipedia.org/wiki/Pope_Clement_XII
Pope Clement XIII	http://en.wikipedia.org/wiki/Pope_Clement_XIII
Pope Clement XIV	http://en.wikipedia.org/wiki/Pope_Clement_XIV
Pope Damasus I	http://en.wikipedia.org/wiki/Pope_Damasus_I
Pope Damasus II	http://en.wikipedia.org/wiki/Pope_Damasus_II
Pope Formosus	http://en.wikipedia.org/wiki/Pope_Formosus
Pope Gregory I	http://en.wikipedia.org/wiki/Pope_Gregory_I
Pope Gregory II	http://en.wikipedia.org/wiki/Pope_Gregory_II
Pope Gregory III	http://en.wikipedia.org/wiki/Pope_Gregory_III
Pope Gregory IV	http://en.wikipedia.org/wiki/Pope_Gregory_IV
Pope Gregory IX	http://en.wikipedia.org/wiki/Pope_Gregory_IX
Pope Gregory V	http://en.wikipedia.org/wiki/Pope_Gregory_V
Pope Gregory VI	http://en.wikipedia.org/wiki/Pope_Gregory_VI
Pope Gregory VII	http://en.wikipedia.org/wiki/Pope_Gregory_VII
Pope Gregory VIII	http://en.wikipedia.org/wiki/Pope_Gregory_VIII
Pope Gregory X	http://en.wikipedia.org/wiki/Pope_Gregory_X
Pope Gregory XI	http://en.wikipedia.org/wiki/Pope_Gregory_XI
Pope Gregory XII	http://en.wikipedia.org/wiki/Pope_Gregory_XII
Pope Gregory XIII	http://en.wikipedia.org/wiki/Pope_Gregory_XIII
Pope Gregory XIV	http://en.wikipedia.org/wiki/Pope_Gregory_XIV
Pope Gregory XV	http://en.wikipedia.org/wiki/Pope_Gregory_XV
Pope Gregory XVI	http://en.wikipedia.org/wiki/Pope_Gregory_XVI
Pope Honorius I	http://en.wikipedia.org/wiki/Pope_Honorius_I
Pope Honorius II	http://en.wikipedia.org/wiki/Pope_Honorius_II
Pope Honorius III	http://en.wikipedia.org/wiki/Pope_Honorius_III
Pope Honorius IV	http://en.wikipedia.org/wiki/Pope_Honorius_IV
Pope Hormisdas	http://en.wikipedia.org/wiki/Pope_Hormisdas
Pope Innocent I	http://en.wikipedia.org/wiki/Pope_Innocent_I
Pope Innocent II	http://en.wikipedia.org/wiki/Pope_Innocent_II
Pope Innocent III	http://en.wikipedia.org/wiki/Pope_Innocent_III
Pope Innocent IV	http://en.wikipedia.org/wiki/Pope_Innocent_IV
Pope Innocent IX	http://en.wikipedia.org/wiki/Pope_Innocent_IX
Pope Innocent V	http://en.wikipedia.org/wiki/Pope_Innocent_V
Pope Innocent VI	http://en.wikipedia.org/wiki/Pope_Innocent_VI
Pope Innocent VII	http://en.wikipedia.org/wiki/Pope_Innocent_VII
Pope Innocent VIII	http://en.wikipedia.org/wiki/Pope_Innocent_VIII
Pope Innocent X	http://en.wikipedia.org/wiki/Pope_Innocent_X
Pope Innocent XI	http://en.wikipedia.org/wiki/Pope_Innocent_XI
Pope Innocent XII	http://en.wikipedia.org/wiki/Pope_Innocent_XII
Pope Innocent XIII	http://en.wikipedia.org/wiki/Pope_Innocent_XIII
Pope John I	http://en.wikipedia.org/wiki/Pope_John_I
Pope John II	http://en.wikipedia.org/wiki/Pope_John_II
Pope John III	http://en.wikipedia.org/wiki/Pope_John_III
Pope John IV	http://en.wikipedia.org/wiki/Pope_John_IV
Pope John IX	http://en.wikipedia.org/wiki/Pope_John_IX
Pope John Paul I	http://en.wikipedia.org/wiki/Pope_John_Paul_I
Pope John Paul II	http://en.wikipedia.org/wiki/Pope_John_Paul_II
Pope John V	http://en.wikipedia.org/wiki/Pope_John_V
Pope John VI	http://en.wikipedia.org/wiki/Pope_John_VI
Pope John VII	http://en.wikipedia.org/wiki/Pope_John_VII
Pope John VIII	http://en.wikipedia.org/wiki/Pope_John_VIII
Pope John X	http://en.wikipedia.org/wiki/Pope_John_X
Pope John XI	http://en.wikipedia.org/wiki/Pope_John_XI
Pope John XII	http://en.wikipedia.org/wiki/Pope_John_XII
Pope John XIII	http://en.wikipedia.org/wiki/Pope_John_XIII
Pope John XIV	http://en.wikipedia.org/wiki/Pope_John_XIV
Pope John XIX	http://en.wikipedia.org/wiki/Pope_John_XIX
Pope John XV	http://en.wikipedia.org/wiki/Pope_John_XV
Pope John XXI	http://en.wikipedia.org/wiki/Pope_John_XXI
Pope John XXII	http://en.wikipedia.org/wiki/Pope_John_XXII
Pope John XXIII	http://en.wikipedia.org/wiki/Pope_John_XXIII
Pope Julius I	http://en.wikipedia.org/wiki/Pope_Julius_I
Pope Julius II	http://en.wikipedia.org/wiki/Pope_Julius_II
Pope Julius III	http://en.wikipedia.org/wiki/Pope_Julius_III
Pope Leo I	http://en.wikipedia.org/wiki/Pope_Leo_I
Pope Leo II	http://en.wikipedia.org/wiki/Pope_Leo_II
Pope Leo III	http://en.wikipedia.org/wiki/Pope_Leo_III
Pope Leo IV	http://en.wikipedia.org/wiki/Pope_Leo_IV
Pope Leo IX	http://en.wikipedia.org/wiki/Pope_Leo_IX
Pope Leo VIII	http://en.wikipedia.org/wiki/Pope_Leo_VIII
Pope Leo X	http://en.wikipedia.org/wiki/Pope_Leo_X
Pope Leo XI	http://en.wikipedia.org/wiki/Pope_Leo_XI
Pope Leo XII	http://en.wikipedia.org/wiki/Pope_Leo_XII
Pope Leo XIII	http://en.wikipedia.org/wiki/Pope_Leo_XIII
Pope Lucius I	http://en.wikipedia.org/wiki/Pope_Lucius_I
Pope Lucius II	http://en.wikipedia.org/wiki/Pope_Lucius_II
Pope Lucius III	http://en.wikipedia.org/wiki/Pope_Lucius_III
Pope Marcellinus	http://en.wikipedia.org/wiki/Pope_Marcellinus
Pope Marcellus I	http://en.wikipedia.org/wiki/Pope_Marcellus_I
Pope Marcellus II	http://en.wikipedia.org/wiki/Pope_Marcellus_II
Pope Marinus I	http://en.wikipedia.org/wiki/Pope_Marinus_I
Pope Marinus II	http://en.wikipedia.org/wiki/Pope_Marinus_II
Pope Nicholas I	http://en.wikipedia.org/wiki/Pope_Nicholas_I
Pope Nicholas II	http://en.wikipedia.org/wiki/Pope_Nicholas_II
Pope Nicholas III	http://en.wikipedia.org/wiki/Pope_Nicholas_III
Pope Paschal I	http://en.wikipedia.org/wiki/Pope_Paschal_I
Pope Paschal II	http://en.wikipedia.org/wiki/Pope_Paschal_II
Pope Paul I	http://en.wikipedia.org/wiki/Pope_Paul_I
Pope Paul II	http://en.wikipedia.org/wiki/Pope_Paul_II
Pope Paul III	http://en.wikipedia.org/wiki/Pope_Paul_III
Pope Paul IV	http://en.wikipedia.org/wiki/Pope_Paul_IV
Pope Paul V	http://en.wikipedia.org/wiki/Pope_Paul_V
Pope Paul VI	http://en.wikipedia.org/wiki/Pope_Paul_VI
Pope Pelagius I	http://en.wikipedia.org/wiki/Pope_Pelagius_I
Pope Pelagius II	http://en.wikipedia.org/wiki/Pope_Pelagius_II
Pope Pius II	http://en.wikipedia.org/wiki/Pope_Pius_II
Pope Pius III	http://en.wikipedia.org/wiki/Pope_Pius_III
Pope Pius IV	http://en.wikipedia.org/wiki/Pope_Pius_IV
Pope Pius IX	http://en.wikipedia.org/wiki/Pope_Pius_IX
Pope Pius V	http://en.wikipedia.org/wiki/Pope_Pius_V
Pope Pius VI	http://en.wikipedia.org/wiki/Pope_Pius_VI
Pope Pius VII	http://en.wikipedia.org/wiki/Pope_Pius_VII
Pope Pius VIII	http://en.wikipedia.org/wiki/Pope_Pius_VIII
Pope Pius X	http://en.wikipedia.org/wiki/Pope_Pius_X
Pope Pius XI	http://en.wikipedia.org/wiki/Pope_Pius_XI
Pope Pius XII	http://en.wikipedia.org/wiki/Pope_Pius_XII
Pope Sergius I	http://en.wikipedia.org/wiki/Pope_Sergius_I
Pope Sergius II	http://en.wikipedia.org/wiki/Pope_Sergius_II
Pope Sergius III	http://en.wikipedia.org/wiki/Pope_Sergius_III
Pope Sixtus III	http://en.wikipedia.org/wiki/Pope_Sixtus_III
Pope Sixtus IV	http://en.wikipedia.org/wiki/Pope_Sixtus_IV
Pope Sixtus V	http://en.wikipedia.org/wiki/Pope_Sixtus_V
Pope Stephen II	http://en.wikipedia.org/wiki/Pope_Stephen_II
Pope Stephen III	http://en.wikipedia.org/wiki/Pope_Stephen_III
Pope Stephen IV	http://en.wikipedia.org/wiki/Pope_Stephen_IV
Pope Stephen IX	http://en.wikipedia.org/wiki/Pope_Stephen_IX
Pope Stephen V	http://en.wikipedia.org/wiki/Pope_Stephen_V
Pope Stephen VI	http://en.wikipedia.org/wiki/Pope_Stephen_VI
Pope Sylvester I	http://en.wikipedia.org/wiki/Pope_Sylvester_I
Pope Symmachus	http://en.wikipedia.org/wiki/Pope_Symmachus
Pope Urban II	http://en.wikipedia.org/wiki/Pope_Urban_II
Pope Urban III	http://en.wikipedia.org/wiki/Pope_Urban_III
Pope Urban IV	http://en.wikipedia.org/wiki/Pope_Urban_IV
Pope Urban V	http://en.wikipedia.org/wiki/Pope_Urban_V
Pope Urban VI	http://en.wikipedia.org/wiki/Pope_Urban_VI
Pope Urban VII	http://en.wikipedia.org/wiki/Pope_Urban_VII
Pope Urban VIII	http://en.wikipedia.org/wiki/Pope_Urban_VIII
Pope Victor I	http://en.wikipedia.org/wiki/Pope_Victor_I
Pope Victor II	http://en.wikipedia.org/wiki/Pope_Victor_II
Pope Victor III	http://en.wikipedia.org/wiki/Pope_Victor_III
Poppy Montgomery	http://en.wikipedia.org/wiki/Poppy_Montgomery
Poppy Z. Brite	http://en.wikipedia.org/wiki/Poppy_Z._Brite
Pops Staples	http://en.wikipedia.org/wiki/Pops_Staples
Porfirio D�az	http://en.wikipedia.org/wiki/Porfirio_D%EDaz
Porfirio Lobo Sosa	http://en.wikipedia.org/wiki/Porfirio_Lobo_Sosa
Porter Goss	http://en.wikipedia.org/wiki/Porter_Goss
Porter Hall	http://en.wikipedia.org/wiki/Porter_Hall
Porter Wagoner	http://en.wikipedia.org/wiki/Porter_Wagoner
Portia de Rossi	http://en.wikipedia.org/wiki/Portia_de_Rossi
Portia Simpson-Miller	http://en.wikipedia.org/wiki/Portia_Simpson-Miller
Potter Stewart	http://en.wikipedia.org/wiki/Potter_Stewart
Poul Anderson	http://en.wikipedia.org/wiki/Poul_Anderson
Poultney Bigelow	http://en.wikipedia.org/wiki/Poultney_Bigelow
Powers Boothe	http://en.wikipedia.org/wiki/Powers_Boothe
Pramoedya Ananta Toer	http://en.wikipedia.org/wiki/Pramoedya_Ananta_Toer
Pratibha Patil	http://en.wikipedia.org/wiki/Pratibha_Patil
Prentiss Ingraham	http://en.wikipedia.org/wiki/Prentiss_Ingraham
Prescott Bush	http://en.wikipedia.org/wiki/Prescott_Bush
Prescott S. Bush, Jr.	http://en.wikipedia.org/wiki/Prescott_S._Bush%2C_Jr.
Preston Sturges	http://en.wikipedia.org/wiki/Preston_Sturges
Primo Levi	http://en.wikipedia.org/wiki/Primo_Levi
Prince Akishino	http://en.wikipedia.org/wiki/Prince_Akishino
Prince Albert II	http://en.wikipedia.org/wiki/Prince_Albert_II
Prince Andrew	http://en.wikipedia.org/wiki/Prince_Andrew
Prince Bandar bin Sultan	http://en.wikipedia.org/wiki/Prince_Bandar_bin_Sultan
Prince Bernhard	http://en.wikipedia.org/wiki/Prince_Bernhard
Prince Buster	http://en.wikipedia.org/wiki/Prince_Buster
Prince Charles	http://en.wikipedia.org/wiki/Prince_Charles
Prince Edward	http://en.wikipedia.org/wiki/Prince_Edward,_Earl_of_Wessex
Prince Ernst August of Hanover	http://en.wikipedia.org/wiki/Prince_Ernst_August_of_Hanover
Prince Frederik	http://en.wikipedia.org/wiki/Prince_Frederik
Prince Hans-Adam II	http://en.wikipedia.org/wiki/Prince_Hans-Adam_II
Prince Harry	http://en.wikipedia.org/wiki/Prince_Harry
Prince Hitachi	http://en.wikipedia.org/wiki/Prince_Hitachi
Prince Lavaka Ata 'Ulukalala	http://en.wikipedia.org/wiki/Prince_Lavaka_Ata_%27Ulukalala
Prince Michael of Kent	http://en.wikipedia.org/wiki/Prince_Michael_of_Kent
Prince Mikasa	http://en.wikipedia.org/wiki/Prince_Mikasa
Prince Naruhito	http://en.wikipedia.org/wiki/Naruhito,_Crown_Prince_of_Japan
Prince of Asturias	http://en.wikipedia.org/wiki/Felipe,_Prince_of_Asturias
Prince Paul	http://en.wikipedia.org/wiki/Prince_Paul_(producer)
Prince Philip	http://en.wikipedia.org/wiki/Prince_Philip
Prince Rainier	http://en.wikipedia.org/wiki/Prince_Rainier
Prince Sultan bin Abdul Aziz	http://en.wikipedia.org/wiki/Prince_Sultan_bin_Abdul_Aziz
Prince William	http://en.wikipedia.org/wiki/Prince_William
Princess Alice	http://en.wikipedia.org/wiki/Princess_Alice,_Duchess_of_Gloucester
Princess Anne	http://en.wikipedia.org/wiki/Princess_Anne
Princess Caroline	http://en.wikipedia.org/wiki/Caroline,_Princess_of_Hanover
Princess Juliana	http://en.wikipedia.org/wiki/Princess_Juliana
Princess Margaret	http://en.wikipedia.org/wiki/Princess_Margaret
Princess Michael of Kent	http://en.wikipedia.org/wiki/Princess_Michael_of_Kent
Princess Stephanie	http://en.wikipedia.org/wiki/Princess_Stéphanie_of_Monaco
Priscilla Barnes	http://en.wikipedia.org/wiki/Priscilla_Barnes
Priscilla Presley	http://en.wikipedia.org/wiki/Priscilla_Presley
Priscilla Taylor	http://en.wikipedia.org/wiki/Priscilla_Taylor
Priti Patel	http://en.wikipedia.org/wiki/Priti_Patel
Professor X	http://en.wikipedia.org/wiki/Professor_X_The_Overseer_(hip_hop)
Prophet Muhammad	http://en.wikipedia.org/wiki/Prophet_Muhammad
Prosper M�rim�e	http://en.wikipedia.org/wiki/Prosper_M%E9rim%E9e
Prospero Alpini	http://en.wikipedia.org/wiki/Prospero_Alpini
Prunella Scales	http://en.wikipedia.org/wiki/Prunella_Scales
Publius Sulpicius Rufus	http://en.wikipedia.org/wiki/Publius_Sulpicius_Rufus
Puff Daddy	http://en.wikipedia.org/wiki/Puff_Daddy
Pyotr Kapitsa	http://en.wikipedia.org/wiki/Pyotr_Kapitsa
Qaboos Bin Said	http://en.wikipedia.org/wiki/Qaboos_Bin_Said
Queen Anne	http://en.wikipedia.org/wiki/Anne_of_Great_Britain
Queen Beatrix I	http://en.wikipedia.org/wiki/Beatrix_of_the_Netherlands
Queen Elizabeth I	http://en.wikipedia.org/wiki/Queen_Elizabeth_I
Queen Elizabeth II	http://en.wikipedia.org/wiki/Queen_Elizabeth_II
Queen Isabella	http://en.wikipedia.org/wiki/Isabella_I_of_Castile
Queen Latifah	http://en.wikipedia.org/wiki/Queen_Latifah
Queen Margrethe II	http://en.wikipedia.org/wiki/Queen_Margrethe_II
Queen Mary I	http://en.wikipedia.org/wiki/Mary_I_of_England
Queen Mary II	http://en.wikipedia.org/wiki/Mary_II_of_England
Queen Noor	http://en.wikipedia.org/wiki/Queen_Noor
Queen Victoria	http://en.wikipedia.org/wiki/Queen_Victoria
Queenie Leonard	http://en.wikipedia.org/wiki/Queenie_Leonard
Quentin Crisp	http://en.wikipedia.org/wiki/Quentin_Crisp
Quentin Kopp	http://en.wikipedia.org/wiki/Quentin_Kopp
Quentin N. Burdick	http://en.wikipedia.org/wiki/Quentin_N._Burdick
Quentin Roosevelt	http://en.wikipedia.org/wiki/Quentin_Roosevelt
Quentin Tarantino	http://en.wikipedia.org/wiki/Quentin_Tarantino
Quincy Jones	http://en.wikipedia.org/wiki/Quincy_Jones
Quinn Martin	http://en.wikipedia.org/wiki/Quinn_Martin
Quintus Ennius	http://en.wikipedia.org/wiki/Quintus_Ennius
Quintus Hortensius	http://en.wikipedia.org/wiki/Quintus_Hortensius
Qusay Hussein	http://en.wikipedia.org/wiki/Qusay_Hussein
R. A. Salvatore	http://en.wikipedia.org/wiki/R._A._Salvatore
R. Buckminster Fuller	http://en.wikipedia.org/wiki/R._Buckminster_Fuller
R. Budd Dwyer	http://en.wikipedia.org/wiki/R._Budd_Dwyer
R. David Paulison	http://en.wikipedia.org/wiki/R._David_Paulison
R. E. Raspe	http://en.wikipedia.org/wiki/R._E._Raspe
R. G. Collingwood	http://en.wikipedia.org/wiki/R._G._Collingwood
R. H. Tawney	http://en.wikipedia.org/wiki/R._H._Tawney
R. J. Rushdoony	http://en.wikipedia.org/wiki/R._J._Rushdoony
R. K. Narayan	http://en.wikipedia.org/wiki/R._K._Narayan
R. Kelly	http://en.wikipedia.org/wiki/R._Kelly
R. L. Burnside	http://en.wikipedia.org/wiki/R._L._Burnside
R. L. Stine	http://en.wikipedia.org/wiki/R._L._Stine
R. Lee Ermey	http://en.wikipedia.org/wiki/R._Lee_Ermey
R. Meredith Belbin	http://en.wikipedia.org/wiki/Meredith_Belbin
R. Michael DeWine	http://en.wikipedia.org/wiki/R._Michael_DeWine
R. Nicholas Burns	http://en.wikipedia.org/wiki/R._Nicholas_Burns
Raab Himself	http://en.wikipedia.org/wiki/Raab_Himself
Rabanus Maurus	http://en.wikipedia.org/wiki/Rabanus_Maurus
Rabih Abou-Khalil	http://en.wikipedia.org/wiki/Rabih_Abou-Khalil
Rabindranath Tagore	http://en.wikipedia.org/wiki/Rabindranath_Tagore
Rachael Leigh Cook	http://en.wikipedia.org/wiki/Rachael_Leigh_Cook
Rachael Ray	http://en.wikipedia.org/wiki/Rachael_Ray
Rachel Bilson	http://en.wikipedia.org/wiki/Rachel_Bilson
Rachel Blanchard	http://en.wikipedia.org/wiki/Rachel_Blanchard
Rachel Carson	http://en.wikipedia.org/wiki/Rachel_Carson
Rachel Corrie	http://en.wikipedia.org/wiki/Rachel_Corrie
Rachel Crothers	http://en.wikipedia.org/wiki/Rachel_Crothers
Rachel Dratch	http://en.wikipedia.org/wiki/Rachel_Dratch
Rachel Griffiths	http://en.wikipedia.org/wiki/Rachel_Griffiths
Rachel Haden	http://en.wikipedia.org/wiki/Rachel_Haden
Rachel Hunter	http://en.wikipedia.org/wiki/Rachel_Hunter
Rachel Kempson	http://en.wikipedia.org/wiki/Rachel_Kempson
Rachel McAdams	http://en.wikipedia.org/wiki/Rachel_McAdams
Rachel Miner	http://en.wikipedia.org/wiki/Rachel_Miner
Rachel Reeves	http://en.wikipedia.org/wiki/Rachel_Reeves
Rachel Shelley	http://en.wikipedia.org/wiki/Rachel_Shelley
Rachel Stevens	http://en.wikipedia.org/wiki/Rachel_Stevens
Rachel Ticotin	http://en.wikipedia.org/wiki/Rachel_Ticotin
Rachel True	http://en.wikipedia.org/wiki/Rachel_True
Rachel Ward	http://en.wikipedia.org/wiki/Rachel_Ward
Rachel Weisz	http://en.wikipedia.org/wiki/Rachel_Weisz
Radha Mitchell	http://en.wikipedia.org/wiki/Radha_Mitchell
Radha Mitchell	http://en.wikipedia.org/wiki/Radha_Mitchell
Radovan Karadzic	http://en.wikipedia.org/wiki/Radovan_Karadzic
Rae Carruth	http://en.wikipedia.org/wiki/Rae_Carruth
Rae Dawn Chong	http://en.wikipedia.org/wiki/Rae_Dawn_Chong
Rafael Alers	http://en.wikipedia.org/wiki/Rafael_Alers
Rafael Alvarez	http://en.wikipedia.org/wiki/Rafael_Alvarez
Rafael Benitez	http://en.wikipedia.org/wiki/Rafael_Benitez
Rafael Correa	http://en.wikipedia.org/wiki/Rafael_Correa
Rafael Le�nidas Trujillo	http://en.wikipedia.org/wiki/Rafael_Le%F3nidas_Trujillo
Rafael Nadal	http://en.wikipedia.org/wiki/Rafael_Nadal
Rafael Palmeiro	http://en.wikipedia.org/wiki/Rafael_Palmeiro
Rafer Johnson	http://en.wikipedia.org/wiki/Rafer_Johnson
Rafik Hariri	http://en.wikipedia.org/wiki/Rafik_Hariri
Ragnar Frisch	http://en.wikipedia.org/wiki/Ragnar_Frisch
Rahm Emanuel	http://en.wikipedia.org/wiki/Rahm_Emanuel
Rahul Dravid	http://en.wikipedia.org/wiki/Rahul_Dravid
Raila Odinga	http://en.wikipedia.org/wiki/Raila_Odinga
Raimondo Montecuccoli	http://en.wikipedia.org/wiki/Raimondo_Montecuccoli
Rainer Barzel	http://en.wikipedia.org/wiki/Rainer_Barzel
Rainer Maria Rilke	http://en.wikipedia.org/wiki/Rainer_Maria_Rilke
Rainer Werner Fassbinder	http://en.wikipedia.org/wiki/Rainer_Werner_Fassbinder
Rainn Wilson	http://en.wikipedia.org/wiki/Rainn_Wilson
Raisa Gorbachev	http://en.wikipedia.org/wiki/Raisa_Gorbachev
Raj Kapoor	http://en.wikipedia.org/wiki/Raj_Kapoor
Rajiv Gandhi	http://en.wikipedia.org/wiki/Rajiv_Gandhi
Ralf H�tter	http://en.wikipedia.org/wiki/Ralf_H%FCtter
Ralph Abercromby	http://en.wikipedia.org/wiki/Ralph_Abercromby
Ralph Abernathy	http://en.wikipedia.org/wiki/Ralph_Abernathy
Ralph Baer	http://en.wikipedia.org/wiki/Ralph_Baer
Ralph Bakshi	http://en.wikipedia.org/wiki/Ralph_Bakshi
Ralph Bellamy	http://en.wikipedia.org/wiki/Ralph_Bellamy
Ralph Bunche	http://en.wikipedia.org/wiki/Ralph_Bunche
Ralph Carter	http://en.wikipedia.org/wiki/Ralph_Carter
Ralph Connor	http://en.wikipedia.org/wiki/Ralph_Connor
Ralph Cooper	http://en.wikipedia.org/wiki/Ralph_Cooper_%28Apollo%29
Ralph Cudworth	http://en.wikipedia.org/wiki/Ralph_Cudworth
Ralph Edwards	http://en.wikipedia.org/wiki/Ralph_Edwards
Ralph Ellison	http://en.wikipedia.org/wiki/Ralph_Ellison
Ralph Fiennes	http://en.wikipedia.org/wiki/Ralph_Fiennes
Ralph Gonsalves	http://en.wikipedia.org/wiki/Ralph_Gonsalves
Ralph Hall	http://en.wikipedia.org/wiki/Ralph_Hall
Ralph Hodgson	http://en.wikipedia.org/wiki/Ralph_Hodgson
Ralph Hopton	http://en.wikipedia.org/wiki/Ralph_Hopton
Ralph Kiner	http://en.wikipedia.org/wiki/Ralph_Kiner
Ralph Lauren	http://en.wikipedia.org/wiki/Ralph_Lauren
Ralph M. Hall	http://en.wikipedia.org/wiki/Ralph_M._Hall
Ralph Macchio	http://en.wikipedia.org/wiki/Ralph_Macchio
Ralph Merkle	http://en.wikipedia.org/wiki/Ralph_Merkle
Ralph Nader	http://en.wikipedia.org/wiki/Ralph_Nader
Ralph Neas	http://en.wikipedia.org/wiki/Ralph_Neas
Ralph Reed	http://en.wikipedia.org/wiki/Ralph_E._Reed,_Jr.
Ralph Regula	http://en.wikipedia.org/wiki/Ralph_Regula
Ralph Richardson	http://en.wikipedia.org/wiki/Ralph_Richardson
Ralph S. Regula	http://en.wikipedia.org/wiki/Ralph_S._Regula
Ralph Sampson	http://en.wikipedia.org/wiki/Ralph_Sampson
Ralph Steadman	http://en.wikipedia.org/wiki/Ralph_Steadman
Ralph Vaughan Williams	http://en.wikipedia.org/wiki/Ralph_Vaughan_Williams
Ralph Waite	http://en.wikipedia.org/wiki/Ralph_Waite
Ralph Waldo Emerson	http://en.wikipedia.org/wiki/Ralph_Waldo_Emerson
Ralph Yarborough	http://en.wikipedia.org/wiki/Ralph_Yarborough
Ram Baran Yadav	http://en.wikipedia.org/wiki/Ram_Baran_Yadav
Ramon Magsaysay	http://en.wikipedia.org/wiki/Ramon_Magsaysay
Ramon Novarro	http://en.wikipedia.org/wiki/Ramon_Novarro
Ramsay MacDonald	http://en.wikipedia.org/wiki/Ramsay_MacDonald
Ramsey Clark	http://en.wikipedia.org/wiki/Ramsey_Clark
Ramzi Yousef	http://en.wikipedia.org/wiki/Ramzi_Yousef
Rand Beers	http://en.wikipedia.org/wiki/Rand_Beers
Randal Cremer	http://en.wikipedia.org/wiki/Randal_Cremer
Randal Kleiser	http://en.wikipedia.org/wiki/Randal_Kleiser
Randall Adams	http://en.wikipedia.org/wiki/Randall_Adams
Randall Jarrell	http://en.wikipedia.org/wiki/Randall_Jarrell
Randall Terry	http://en.wikipedia.org/wiki/Randall_Terry
Randi Rhodes	http://en.wikipedia.org/wiki/Randi_Rhodes
Randolph Churchill	http://en.wikipedia.org/wiki/Randolph_Churchill
Randolph Mantooth	http://en.wikipedia.org/wiki/Randolph_Mantooth
Randolph Scott	http://en.wikipedia.org/wiki/Randolph_Scott
Randy Bachman	http://en.wikipedia.org/wiki/Randy_Bachman
Randy Castillo	http://en.wikipedia.org/wiki/Randy_Castillo
Randy DeBarge	http://en.wikipedia.org/wiki/Randy_DeBarge
Randy Forbes	http://en.wikipedia.org/wiki/Randy_Forbes
Randy Gardner	http://en.wikipedia.org/wiki/Randy_Gardner_(figure_skater)
Randy Harrison	http://en.wikipedia.org/wiki/Randy_Harrison
Randy Jackson	http://en.wikipedia.org/wiki/Randy_Jackson
Randy Johnson	http://en.wikipedia.org/wiki/Randy_Johnson
Randy Kuhl	http://en.wikipedia.org/wiki/Randy_Kuhl
Randy Moss	http://en.wikipedia.org/wiki/Randy_Moss
Randy Neugebauer	http://en.wikipedia.org/wiki/Randy_Neugebauer
Randy Newman	http://en.wikipedia.org/wiki/Randy_Newman
Randy Orton	http://en.wikipedia.org/wiki/Randy_Orton
Randy Quaid	http://en.wikipedia.org/wiki/Randy_Quaid
Randy Rhoads	http://en.wikipedia.org/wiki/Randy_Rhoads
Randy Savage	http://en.wikipedia.org/wiki/Randy_Savage
Randy Travis	http://en.wikipedia.org/wiki/Randy_Travis
Randy Warmer	http://en.wikipedia.org/wiki/Randy_VanWarmer
Randy Weaver	http://en.wikipedia.org/wiki/Randy_Weaver
Raoul Dufy	http://en.wikipedia.org/wiki/Raoul_Dufy
Raoul Wallenberg	http://en.wikipedia.org/wiki/Raoul_Wallenberg
Raoul Walsh	http://en.wikipedia.org/wiki/Raoul_Walsh
Raphael Holinshed	http://en.wikipedia.org/wiki/Raphael_Holinshed
Raphael Saadiq	http://en.wikipedia.org/wiki/Raphael_Saadiq
Raquel Alessi	http://en.wikipedia.org/wiki/Raquel_Alessi
Raquel Welch	http://en.wikipedia.org/wiki/Raquel_Welch
Rasheed Wallace	http://en.wikipedia.org/wiki/Rasheed_Wallace
Rashid Khalidi	http://en.wikipedia.org/wiki/Rashid_Khalidi
Rashida Jones	http://en.wikipedia.org/wiki/Rashida_Jones
Rasmus B. Anderson	http://en.wikipedia.org/wiki/Rasmus_B._Anderson
Ratnasiri Wickremanayake	http://en.wikipedia.org/wiki/Ratnasiri_Wickremanayake
Ratu Josefa Iloilo	http://en.wikipedia.org/wiki/Ratu_Josefa_Iloilo
Ra�l Alfons�n	http://en.wikipedia.org/wiki/Ra%FAl_Alfons%EDn
Ra�l Castro	http://en.wikipedia.org/wiki/Ra%FAl_Castro
Ra�l Grijalva	http://en.wikipedia.org/wiki/Ra%FAl_Grijalva
Raul Julia	http://en.wikipedia.org/wiki/Raul_Julia
Ravi Shankar	http://en.wikipedia.org/wiki/Ravi_Shankar
Ray Anthony	http://en.wikipedia.org/wiki/Ray_Anthony
Ray Benzino	http://en.wikipedia.org/wiki/Ray_Benzino
Ray Bolger	http://en.wikipedia.org/wiki/Ray_Bolger
Ray Bradbury	http://en.wikipedia.org/wiki/Ray_Bradbury
Ray Charles	http://en.wikipedia.org/wiki/Ray_Charles
Ray Collins	http://en.wikipedia.org/wiki/Ray_Collins_(actor)
Ray Combs	http://en.wikipedia.org/wiki/Ray_Combs
Ray Davies	http://en.wikipedia.org/wiki/Ray_Davies
Ray Goulding	http://en.wikipedia.org/wiki/Ray_Goulding
Ray Harryhausen	http://en.wikipedia.org/wiki/Ray_Harryhausen
Ray Kroc	http://en.wikipedia.org/wiki/Ray_Kroc
Ray Kurzweil	http://en.wikipedia.org/wiki/Ray_Kurzweil
Ray LaHood	http://en.wikipedia.org/wiki/Ray_LaHood
Ray Lewis	http://en.wikipedia.org/wiki/Ray_Lewis
Ray Liotta	http://en.wikipedia.org/wiki/Ray_Liotta
Ray Manzarek	http://en.wikipedia.org/wiki/Ray_Manzarek
Ray Marshall	http://en.wikipedia.org/wiki/Ray_Marshall
Ray Milland	http://en.wikipedia.org/wiki/Ray_Milland
Ray Nagin	http://en.wikipedia.org/wiki/Ray_Nagin
Ray Noorda	http://en.wikipedia.org/wiki/Ray_Noorda
Ray Price	http://en.wikipedia.org/wiki/Ray_Price_(musician)
Ray Romano	http://en.wikipedia.org/wiki/Ray_Romano
Ray Sharkey	http://en.wikipedia.org/wiki/Ray_Sharkey
Ray Stannard Baker	http://en.wikipedia.org/wiki/Ray_Stannard_Baker
Ray Stevens	http://en.wikipedia.org/wiki/Ray_Stevens
Ray Suarez	http://en.wikipedia.org/wiki/Ray_Suarez
Ray Taliaferro	http://en.wikipedia.org/wiki/Ray_Taliaferro
Ray Toro	http://en.wikipedia.org/wiki/Ray_Toro
Ray Walston	http://en.wikipedia.org/wiki/Ray_Walston
Ray Wise	http://en.wikipedia.org/wiki/Ray_Wise
Raymond A. Hare	http://en.wikipedia.org/wiki/Raymond_A._Hare
Raymond Bailey	http://en.wikipedia.org/wiki/Raymond_Bailey
Raymond Barre	http://en.wikipedia.org/wiki/Raymond_Barre
Raymond Burr	http://en.wikipedia.org/wiki/Raymond_Burr
Raymond Carver	http://en.wikipedia.org/wiki/Raymond_Carver
Raymond Chandler	http://en.wikipedia.org/wiki/Raymond_Chandler
Raymond Davis, Jr.	http://en.wikipedia.org/wiki/Raymond_Davis%2C_Jr.
Raymond E. Feist	http://en.wikipedia.org/wiki/Raymond_E._Feist
Raymond J. Donovan	http://en.wikipedia.org/wiki/Raymond_J._Donovan
Raymond J. McGrath	http://en.wikipedia.org/wiki/Raymond_J._McGrath
Raymond Lull	http://en.wikipedia.org/wiki/Raymond_Lull
Raymond Massey	http://en.wikipedia.org/wiki/Raymond_Massey
Raymond P. Kogovsek	http://en.wikipedia.org/wiki/Raymond_P._Kogovsek
Raymond Queneau	http://en.wikipedia.org/wiki/Raymond_Queneau
Raymond Radiguet	http://en.wikipedia.org/wiki/Raymond_Radiguet
Raymond Rubicam	http://en.wikipedia.org/wiki/Raymond_Rubicam
Raymond Scott	http://en.wikipedia.org/wiki/Raymond_Scott
Raymond Williams	http://en.wikipedia.org/wiki/Raymond_Williams
Razaaq Adoti	http://en.wikipedia.org/wiki/Razaaq_Adoti
Reba McEntire	http://en.wikipedia.org/wiki/Reba_McEntire
Rebecca De Mornay	http://en.wikipedia.org/wiki/Rebecca_De_Mornay
Rebecca Gayheart	http://en.wikipedia.org/wiki/Rebecca_Gayheart
Rebecca Hagelin	http://en.wikipedia.org/wiki/Rebecca_Hagelin
Rebecca Harris	http://en.wikipedia.org/wiki/Rebecca_Harris
Rebecca Latimer Felton	http://en.wikipedia.org/wiki/Rebecca_Latimer_Felton
Rebecca Loos	http://en.wikipedia.org/wiki/Rebecca_Loos
Rebecca Romijn	http://en.wikipedia.org/wiki/Rebecca_Romijn
Rebecca West	http://en.wikipedia.org/wiki/Rebecca_West
Recep Tayyip Erdogan	http://en.wikipedia.org/wiki/Recep_Tayyip_Erdogan
Red Adair	http://en.wikipedia.org/wiki/Red_Adair
Red Auerbach	http://en.wikipedia.org/wiki/Red_Auerbach
Red Barber	http://en.wikipedia.org/wiki/Red_Barber
Red Buttons	http://en.wikipedia.org/wiki/Red_Buttons
Red Foley	http://en.wikipedia.org/wiki/Red_Foley
Red Skelton	http://en.wikipedia.org/wiki/Red_Skelton
Red Sovine	http://en.wikipedia.org/wiki/Red_Sovine
Redd Foxx	http://en.wikipedia.org/wiki/Redd_Foxx
Reed E. Hundt	http://en.wikipedia.org/wiki/Reed_E._Hundt
Reed Hadley	http://en.wikipedia.org/wiki/Reed_Hadley
Reed Whittemore	http://en.wikipedia.org/wiki/Reed_Whittemore
Reese Witherspoon	http://en.wikipedia.org/wiki/Reese_Witherspoon
Reeves Gabrels	http://en.wikipedia.org/wiki/Reeves_Gabrels
Reg Varney	http://en.wikipedia.org/wiki/Reg_Varney
Reggie Bush	http://en.wikipedia.org/wiki/Reggie_Bush
Reggie Jackson	http://en.wikipedia.org/wiki/Reggie_Jackson
Reggie Miller	http://en.wikipedia.org/wiki/Reggie_Miller
Reggie White	http://en.wikipedia.org/wiki/Reggie_White
Regimantas Adomaitis	http://en.wikipedia.org/wiki/Regimantas_Adomaitis
Regina Hall	http://en.wikipedia.org/wiki/Regina_Hall
Regina King	http://en.wikipedia.org/wiki/Regina_King
Regina M. Anderson	http://en.wikipedia.org/wiki/Regina_M._Anderson
Reginald Denny	http://en.wikipedia.org/wiki/Reginald_Denny_incident
Reginald Denny	http://en.wikipedia.org/wiki/Reginald_Denny_(actor)
Reginald Marsh	http://en.wikipedia.org/wiki/Reginald_Marsh_(artist)
Reginald Owen	http://en.wikipedia.org/wiki/Reginald_Owen
Reginald Punnett	http://en.wikipedia.org/wiki/Reginald_Punnett
Reginald VelJohnson	http://en.wikipedia.org/wiki/Reginald_VelJohnson
Regis Philbin	http://en.wikipedia.org/wiki/Regis_Philbin
Regis Toomey	http://en.wikipedia.org/wiki/Regis_Toomey
Rehman Chishti	http://en.wikipedia.org/wiki/Rehman_Chishti
Reinaldo Arenas	http://en.wikipedia.org/wiki/Reinaldo_Arenas
Reinhard Bonnke	http://en.wikipedia.org/wiki/Reinhard_Bonnke
Reinhard Hardegen	http://en.wikipedia.org/wiki/Reinhard_Hardegen
Reinhard Heydrich	http://en.wikipedia.org/wiki/Reinhard_Heydrich
Reinhold Niebuhr	http://en.wikipedia.org/wiki/Reinhold_Niebuhr
R�my de Gourmont	http://en.wikipedia.org/wiki/R%E9my_de_Gourmont
Rena Sofer	http://en.wikipedia.org/wiki/Rena_Sofer
Renata Adler	http://en.wikipedia.org/wiki/Renata_Adler
Ren� Auberjonois	http://en.wikipedia.org/wiki/René_Auberjonois_(actor)
Ren� Cailli�	http://en.wikipedia.org/wiki/Ren%E9_Cailli%E9
Ren� Cassin	http://en.wikipedia.org/wiki/Ren%E9_Cassin
Ren� Clair	http://en.wikipedia.org/wiki/Ren%E9_Clair
Ren� Descartes	http://en.wikipedia.org/wiki/Ren%E9_Descartes
Ren� L�vesque	http://en.wikipedia.org/wiki/Ren%E9_L%E9vesque
R�n� Louiche Desfontaines	http://en.wikipedia.org/wiki/Ren%C3%A9_Louiche_Desfontaines
Ren� Magritte	http://en.wikipedia.org/wiki/Ren%E9_Magritte
Ren� Marqu�s	http://en.wikipedia.org/wiki/Ren%E9_Marqu%E9s
Ren� Pr�val	http://en.wikipedia.org/wiki/Ren%E9_Pr%E9val
Rene Rivkin	http://en.wikipedia.org/wiki/Rene_Rivkin
Rene Russo	http://en.wikipedia.org/wiki/Rene_Russo
Ren�-Antoine Ferchault de R�aumur	http://en.wikipedia.org/wiki/Ren%E9-Antoine_Ferchault_de_R%E9aumur
Ren�e Ador�e	http://en.wikipedia.org/wiki/Ren%E9e_Ador%E9e
Ren�e O'Connor	http://en.wikipedia.org/wiki/Ren%E9e_O%27Connor
Ren�e Taylor	http://en.wikipedia.org/wiki/Ren%E9e_Taylor
Ren�e Zellweger	http://en.wikipedia.org/wiki/Ren%E9e_Zellweger
Ren�-Just Ha�y	http://en.wikipedia.org/wiki/Ren%E9-Just_Ha%FCy
Renny Harlin	http://en.wikipedia.org/wiki/Renny_Harlin
Renzo Piano	http://en.wikipedia.org/wiki/Renzo_Piano
Retief Goosen	http://en.wikipedia.org/wiki/Retief_Goosen
Reto Salimbeni	http://en.wikipedia.org/wiki/Reto_Salimbeni
Reubin Askew	http://en.wikipedia.org/wiki/Reubin_Askew
Rev. Cecil Williams	http://en.wikipedia.org/wiki/Cecil_Williams
Reverdy Johnson	http://en.wikipedia.org/wiki/Reverdy_Johnson
Rex Allen	http://en.wikipedia.org/wiki/Rex_Allen
Rex Brown	http://en.wikipedia.org/wiki/Rex_Brown
Rex Harrison	http://en.wikipedia.org/wiki/Rex_Harrison
Rex Humbard	http://en.wikipedia.org/wiki/Rex_Humbard
Rex Reed	http://en.wikipedia.org/wiki/Rex_Reed
Rex Stout	http://en.wikipedia.org/wiki/Rex_Stout
Reynolds Price	http://en.wikipedia.org/wiki/Reynolds_Price
Rhea Perlman	http://en.wikipedia.org/wiki/Rhea_Perlman
Rhodri Morgan	http://en.wikipedia.org/wiki/Rhodri_Morgan
Rhona Mitra	http://en.wikipedia.org/wiki/Rhona_Mitra
Rhonda Fleming	http://en.wikipedia.org/wiki/Rhonda_Fleming
Rhys Ifans	http://en.wikipedia.org/wiki/Rhys_Ifans
Ric Flair	http://en.wikipedia.org/wiki/Ric_Flair
Ric Keller	http://en.wikipedia.org/wiki/Ric_Keller
Ric Ocasek	http://en.wikipedia.org/wiki/Ric_Ocasek
Ricardo Flores Mag�n	http://en.wikipedia.org/wiki/Ricardo_Flores_Mag%F3n
Ricardo Franco	http://en.wikipedia.org/wiki/Ricardo_Franco
Ricardo Lagos	http://en.wikipedia.org/wiki/Ricardo_Lagos
Ricardo Lagos	http://en.wikipedia.org/wiki/Ricardo_Lagos
Ricardo Maduro	http://en.wikipedia.org/wiki/Ricardo_Maduro
Ricardo Martinelli	http://en.wikipedia.org/wiki/Ricardo_Martinelli
Ricardo Montalban	http://en.wikipedia.org/wiki/Ricardo_Montalban
Ricardo Piglia	http://en.wikipedia.org/wiki/Ricardo_Piglia
Ricardo Sanchez	http://en.wikipedia.org/wiki/Ricardo_Sanchez
Riccardo Giacconi	http://en.wikipedia.org/wiki/Riccardo_Giacconi
Rich Galen	http://en.wikipedia.org/wiki/Rich_Galen
Rich Hall	http://en.wikipedia.org/wiki/Rich_Hall
Rich Little	http://en.wikipedia.org/wiki/Rich_Little
Rich Lowry	http://en.wikipedia.org/wiki/Rich_Lowry
Rich Robinson	http://en.wikipedia.org/wiki/Rich_Robinson
Richard A. Clarke	http://en.wikipedia.org/wiki/Richard_A._Clarke
Richard A. Gephardt	http://en.wikipedia.org/wiki/Richard_A._Gephardt
Richard Adams	http://en.wikipedia.org/wiki/Richard_Adams
Richard Albrecht	http://en.wikipedia.org/wiki/Richard_Albrecht
Richard Allen	http://en.wikipedia.org/wiki/Richard_Allen_(bishop)
Richard Allen Davis	http://en.wikipedia.org/wiki/Richard_Allen_Davis
Richard Anderson	http://en.wikipedia.org/wiki/Richard_Anderson
Richard Arlen	http://en.wikipedia.org/wiki/Richard_Arlen
Richard Armitage	http://en.wikipedia.org/wiki/Richard_Armitage_(politician)
Richard Ashcroft	http://en.wikipedia.org/wiki/Richard_Ashcroft
Richard Attenborough	http://en.wikipedia.org/wiki/Richard_Attenborough
Richard Avedon	http://en.wikipedia.org/wiki/Richard_Avedon
Richard Ayoade	http://en.wikipedia.org/wiki/Richard_Ayoade
Richard B. Russell	http://en.wikipedia.org/wiki/Richard_Russell,_Jr.
Richard Bach	http://en.wikipedia.org/wiki/Richard_Bach
Richard Bacon	http://en.wikipedia.org/wiki/Richard_Bacon_(politician)
Richard Baker	http://en.wikipedia.org/wiki/Richard_Baker_(U.S._politician)
Richard Barthelmess	http://en.wikipedia.org/wiki/Richard_Barthelmess
Richard Basehart	http://en.wikipedia.org/wiki/Richard_Basehart
Richard Bedford Bennett	http://en.wikipedia.org/wiki/Richard_Bedford_Bennett
Richard Belzer	http://en.wikipedia.org/wiki/Richard_Belzer
Richard Benjamin	http://en.wikipedia.org/wiki/Richard_Benjamin
Richard Bentley	http://en.wikipedia.org/wiki/Richard_Bentley
Richard Ben-Veniste	http://en.wikipedia.org/wiki/Richard_Ben-Veniste
Richard Benyon	http://en.wikipedia.org/wiki/Richard_Benyon
Richard Berry	http://en.wikipedia.org/wiki/Richard_Berry
Richard Beymer	http://en.wikipedia.org/wiki/Richard_Beymer
Richard Biggs	http://en.wikipedia.org/wiki/Richard_Biggs
Richard Boone	http://en.wikipedia.org/wiki/Richard_Boone
Richard Branson	http://en.wikipedia.org/wiki/Richard_Branson
Richard Brautigan	http://en.wikipedia.org/wiki/Richard_Brautigan
Richard Briers	http://en.wikipedia.org/wiki/Richard_Briers
Richard Brinsley Sheridan	http://en.wikipedia.org/wiki/Richard_Brinsley_Sheridan
Richard Brooks	http://en.wikipedia.org/wiki/Richard_Brooks
Richard Bryan	http://en.wikipedia.org/wiki/Richard_Bryan
Richard Burden	http://en.wikipedia.org/wiki/Richard_Burden
Richard Burdon Haldane	http://en.wikipedia.org/wiki/Richard_Burdon_Haldane
Richard Burr	http://en.wikipedia.org/wiki/Richard_Burr
Richard Burton	http://en.wikipedia.org/wiki/Richard_Burton
Richard C. Holbrooke	http://en.wikipedia.org/wiki/Richard_C._Holbrooke
Richard C. Levin	http://en.wikipedia.org/wiki/Richard_C._Levin
Richard C. Notebaert	http://en.wikipedia.org/wiki/Richard_Notebaert
Richard C. Shelby	http://en.wikipedia.org/wiki/Richard_C._Shelby
Richard Carpenter	http://en.wikipedia.org/wiki/Richard_Carpenter_(musician)
Richard Chamberlain	http://en.wikipedia.org/wiki/Richard_Chamberlain
Richard Crenna	http://en.wikipedia.org/wiki/Richard_Crenna
Richard Cromwell	http://en.wikipedia.org/wiki/Richard_Cromwell
Richard D. Fairbank	http://en.wikipedia.org/wiki/Richard_D._Fairbank
Richard D. James	http://en.wikipedia.org/wiki/Richard_D._James
Richard Darman	http://en.wikipedia.org/wiki/Richard_Darman
Richard Dawes	http://en.wikipedia.org/wiki/Richard_Dawes
Richard Dawkins	http://en.wikipedia.org/wiki/Richard_Dawkins
Richard Dawson	http://en.wikipedia.org/wiki/Richard_Dawson
Richard de Bury	http://en.wikipedia.org/wiki/Richard_de_Bury
Richard Deacon	http://en.wikipedia.org/wiki/Richard_Deacon_(actor)
Richard Dean Anderson	http://en.wikipedia.org/wiki/Richard_Dean_Anderson
Richard Deane	http://en.wikipedia.org/wiki/Richard_Deane
Richard Dedekind	http://en.wikipedia.org/wiki/Richard_Dedekind
Richard Denning	http://en.wikipedia.org/wiki/Richard_Denning
Richard Donner	http://en.wikipedia.org/wiki/Richard_Donner
Richard Dorfmeister	http://en.wikipedia.org/wiki/Richard_Dorfmeister
Richard Drax	http://en.wikipedia.org/wiki/Richard_Drax
Richard Dreyfuss	http://en.wikipedia.org/wiki/Richard_Dreyfuss
Richard Durbin	http://en.wikipedia.org/wiki/Dick_Durbin
Richard E. Byrd	http://en.wikipedia.org/wiki/Richard_E._Byrd
Richard E. Grant	http://en.wikipedia.org/wiki/Richard_E._Grant
Richard E. Smalley	http://en.wikipedia.org/wiki/Richard_E._Smalley
Richard E. Taylor	http://en.wikipedia.org/wiki/Richard_E._Taylor
Richard Eberhart	http://en.wikipedia.org/wiki/Richard_Eberhart
Richard Egan	http://en.wikipedia.org/wiki/Richard_Egan_(actor)
Richard Elfman	http://en.wikipedia.org/wiki/Richard_Elfman
Richard Epstein	http://en.wikipedia.org/wiki/Richard_Epstein
Richard F. Outcault	http://en.wikipedia.org/wiki/Richard_F._Outcault
Richard Fanshawe	http://en.wikipedia.org/wiki/Sir_Richard_Fanshawe,_1st_Baronet
Richard Farnsworth	http://en.wikipedia.org/wiki/Richard_Farnsworth
Richard Fell	http://en.wikipedia.org/wiki/Richard_Fell
Richard Feynman	http://en.wikipedia.org/wiki/Richard_Feynman
Richard Fleischer	http://en.wikipedia.org/wiki/Richard_Fleischer
Richard Ford	http://en.wikipedia.org/wiki/Richard_Ford
Richard Fuller	http://en.wikipedia.org/wiki/Richard_Fuller_(politician)
Richard G. Butler	http://en.wikipedia.org/wiki/Richard_G._Butler
Richard G. Lugar	http://en.wikipedia.org/wiki/Richard_G._Lugar
Richard G. Stern	http://en.wikipedia.org/wiki/Richard_G._Stern
Richard Gere	http://en.wikipedia.org/wiki/Richard_Gere
Richard Graham	http://en.wikipedia.org/wiki/Richard_Graham_(politician)
Richard Grasso	http://en.wikipedia.org/wiki/Richard_Grasso
Richard Grieco	http://en.wikipedia.org/wiki/Richard_Grieco
Richard H. Anderson	http://en.wikipedia.org/wiki/Richard_H._Anderson
Richard H. Carmona	http://en.wikipedia.org/wiki/Richard_H._Carmona
Richard H. Lehman	http://en.wikipedia.org/wiki/Richard_H._Lehman
Richard Hakluyt	http://en.wikipedia.org/wiki/Richard_Hakluyt
Richard Harding Davis	http://en.wikipedia.org/wiki/Richard_Harding_Davis
Richard Harrington	http://en.wikipedia.org/wiki/Richard_Harrington_(British_politician)
Richard Harris	http://en.wikipedia.org/wiki/Richard_Harris
Richard Hatch	http://en.wikipedia.org/wiki/Richard_Hatch
Richard Hatch	http://en.wikipedia.org/wiki/Richard_Hatch_(Survivor_contestant)
Richard Haydn	http://en.wikipedia.org/wiki/Richard_Haydn
Richard Hell	http://en.wikipedia.org/wiki/Richard_Hell
Richard Helms	http://en.wikipedia.org/wiki/Richard_Helms
Richard Henry Dana	http://en.wikipedia.org/wiki/Richard_Henry_Dana,_Jr.
Richard Henry Lee	http://en.wikipedia.org/wiki/Richard_Henry_Lee
Richard Henry Stoddard	http://en.wikipedia.org/wiki/Richard_Henry_Stoddard
Richard Hofstadter	http://en.wikipedia.org/wiki/Richard_Hofstadter
Richard Hooker	http://en.wikipedia.org/wiki/Richard_Hooker
Richard Howard	http://en.wikipedia.org/wiki/Richard_Howard
Richard Howe	http://en.wikipedia.org/wiki/Richard_Howe
Richard Hughes	http://en.wikipedia.org/wiki/Richard_Hughes_(writer)
Richard J. Codey	http://en.wikipedia.org/wiki/Richard_J._Codey
Richard J. Daley	http://en.wikipedia.org/wiki/Richard_J._Daley
Richard J. Durbin	http://en.wikipedia.org/wiki/Richard_J._Durbin
Richard Jago	http://en.wikipedia.org/wiki/Richard_Jago
Richard Jewell	http://en.wikipedia.org/wiki/Richard_Jewell
Richard Johnson	http://en.wikipedia.org/wiki/Richard_Johnson_(actor)
Richard Jordan	http://en.wikipedia.org/wiki/Richard_Jordan
Richard Jordan Gatling	http://en.wikipedia.org/wiki/Richard_Jordan_Gatling
Richard K. Armey	http://en.wikipedia.org/wiki/Richard_K._Armey
Richard Karn	http://en.wikipedia.org/wiki/Richard_Karn
Richard Kelly	http://en.wikipedia.org/wiki/Richard_Kelly_(director)
Richard Kelly	http://en.wikipedia.org/wiki/Richard_Kelly_(politician)
Richard Kern	http://en.wikipedia.org/wiki/Richard_Kern
Richard Kiel	http://en.wikipedia.org/wiki/Richard_Kiel
Richard Kiley	http://en.wikipedia.org/wiki/Richard_Kiley
Richard Kirk	http://en.wikipedia.org/wiki/Richard_H._Kirk
Richard Kline	http://en.wikipedia.org/wiki/Richard_Kline
Richard Kostelanetz	http://en.wikipedia.org/wiki/Richard_Kostelanetz
Richard Kuhn	http://en.wikipedia.org/wiki/Richard_Kuhn
Richard L. M. Synge	http://en.wikipedia.org/wiki/Richard_Laurence_Millington_Synge
Richard Land	http://en.wikipedia.org/wiki/Richard_Land
Richard Leakey	http://en.wikipedia.org/wiki/Richard_Leakey
Richard Lepsius	http://en.wikipedia.org/wiki/Richard_Lepsius
Richard Lester	http://en.wikipedia.org/wiki/Richard_Lester
Richard Lewis	http://en.wikipedia.org/wiki/Richard_Lewis_(comedian)
Richard Linklater	http://en.wikipedia.org/wiki/Richard_Linklater
Richard Llewellyn	http://en.wikipedia.org/wiki/Richard_Llewellyn
Richard Long	http://en.wikipedia.org/wiki/Richard_Long_(actor)
Richard Lovelace	http://en.wikipedia.org/wiki/Richard_Lovelace
Richard M. Daley	http://en.wikipedia.org/wiki/Richard_M._Daley
Richard M. Kovacevich	http://en.wikipedia.org/wiki/Richard_Kovacevich
Richard M. Nixon	http://en.wikipedia.org/wiki/Richard_M._Nixon
Richard Manuel	http://en.wikipedia.org/wiki/Richard_Manuel
Richard Marx	http://en.wikipedia.org/wiki/Richard_Marx
Richard Masur	http://en.wikipedia.org/wiki/Richard_Masur
Richard Mentor Johnson	http://en.wikipedia.org/wiki/Richard_Mentor_Johnson
Richard Moll	http://en.wikipedia.org/wiki/Richard_Moll
Richard Monckton Milnes	http://en.wikipedia.org/wiki/Richard_Monckton_Milnes
Richard Montgomery	http://en.wikipedia.org/wiki/Richard_Montgomery
Richard Mulligan	http://en.wikipedia.org/wiki/Richard_Mulligan
Richard Myers	http://en.wikipedia.org/wiki/Richard_Myers
Richard Neal	http://en.wikipedia.org/wiki/Richard_Neal
Richard Neville	http://en.wikipedia.org/wiki/Richard_Neville,_16th_Earl_of_Warwick
Richard Norman Shaw	http://en.wikipedia.org/wiki/Richard_Norman_Shaw
Richard Nugent	http://en.wikipedia.org/wiki/Richard_Bruce_Nugent
Richard O'Brien	http://en.wikipedia.org/wiki/Richard_O%27Brien
Richard Olney	http://en.wikipedia.org/wiki/Richard_Olney
Richard Ottaway	http://en.wikipedia.org/wiki/Richard_Ottaway
Richard Parsons	http://en.wikipedia.org/wiki/Richard_Parsons_(businessman)
Richard Paul	http://en.wikipedia.org/wiki/Richard_Paul
Richard Perle	http://en.wikipedia.org/wiki/Richard_Perle
Richard Petty	http://en.wikipedia.org/wiki/Richard_Petty
Richard Pini	http://en.wikipedia.org/wiki/Richard_Pini
Richard Pombo	http://en.wikipedia.org/wiki/Richard_Pombo
Richard Powers	http://en.wikipedia.org/wiki/Richard_Powers
Richard Pryor	http://en.wikipedia.org/wiki/Richard_Pryor
Richard R. Ernst	http://en.wikipedia.org/wiki/Richard_R._Ernst
Richard Ramirez	http://en.wikipedia.org/wiki/Richard_Ramirez
Richard Ray	http://en.wikipedia.org/wiki/Richard_Ray
Richard Reid	http://en.wikipedia.org/wiki/Richard_Reid_(shoe_bomber)
Richard Rodgers	http://en.wikipedia.org/wiki/Richard_Rodgers
Richard Rodriguez	http://en.wikipedia.org/wiki/Richard_Rodriguez
Richard Roeper	http://en.wikipedia.org/wiki/Richard_Roeper
Richard Rogers	http://en.wikipedia.org/wiki/Richard_Rogers
Richard Rorty	http://en.wikipedia.org/wiki/Richard_Rorty
Richard Roundtree	http://en.wikipedia.org/wiki/Richard_Roundtree
Richard Ruccolo	http://en.wikipedia.org/wiki/Richard_Ruccolo
Richard Rush	http://en.wikipedia.org/wiki/Richard_Rush
Richard Russo	http://en.wikipedia.org/wiki/Richard_Russo
Richard S. Castellano	http://en.wikipedia.org/wiki/Richard_S._Castellano
Richard S. Fuld Jr.	http://en.wikipedia.org/wiki/Richard_S._Fuld_Jr.
Richard Sanders	http://en.wikipedia.org/wiki/Richard_Sanders_(actor)
Richard Savage	http://en.wikipedia.org/wiki/Richard_Savage
Richard Scaife	http://en.wikipedia.org/wiki/Richard_Scaife
Richard Scarry	http://en.wikipedia.org/wiki/Richard_Scarry
Richard Schiff	http://en.wikipedia.org/wiki/Richard_Schiff
Richard Scrushy	http://en.wikipedia.org/wiki/Richard_Scrushy
Richard Shelby	http://en.wikipedia.org/wiki/Richard_Shelby
Richard Shepherd	http://en.wikipedia.org/wiki/Richard_Shepherd
Richard Simmons	http://en.wikipedia.org/wiki/Richard_Simmons
Richard Sorge	http://en.wikipedia.org/wiki/Richard_Sorge
Richard Speck	http://en.wikipedia.org/wiki/Richard_Speck
Richard Stallings	http://en.wikipedia.org/wiki/Richard_Stallings
Richard Stallman	http://en.wikipedia.org/wiki/Richard_Stallman
Richard Steele	http://en.wikipedia.org/wiki/Richard_Steele
Richard Stengel	http://en.wikipedia.org/wiki/Richard_Stengel
Richard Stone	http://en.wikipedia.org/wiki/Richard_Stone
Richard Strauss	http://en.wikipedia.org/wiki/Richard_Strauss
Richard T. Ely	http://en.wikipedia.org/wiki/Richard_T._Ely
Richard Thomas	http://en.wikipedia.org/wiki/Richard_Thomas_(actor)
Richard Thompson	http://en.wikipedia.org/wiki/Richard_Thompson_(musician)
Richard Thorpe	http://en.wikipedia.org/wiki/Richard_Thorpe
Richard Todd	http://en.wikipedia.org/wiki/Richard_Todd
Richard Trethewey	http://en.wikipedia.org/wiki/Richard_Trethewey
Richard V. Allen	http://en.wikipedia.org/wiki/Richard_V._Allen
Richard von Weizs�cker	http://en.wikipedia.org/wiki/Richard_von_Weizs%E4cker
Richard W. Riley	http://en.wikipedia.org/wiki/Richard_W._Riley
Richard W. Sears	http://en.wikipedia.org/wiki/Richard_W._Sears
Richard Wagner	http://en.wikipedia.org/wiki/Richard_Wagner
Richard Widmark	http://en.wikipedia.org/wiki/Richard_Widmark
Richard Wilbur	http://en.wikipedia.org/wiki/Richard_Wilbur
Richard Willst�tter	http://en.wikipedia.org/wiki/Richard_Willst%E4tter
Richard Wright	http://en.wikipedia.org/wiki/Richard_Wright_(author)
Richard Zsigmondy	http://en.wikipedia.org/wiki/Richard_Zsigmondy
Richie Sambora	http://en.wikipedia.org/wiki/Richie_Sambora
Richmond Lattimore	http://en.wikipedia.org/wiki/Richmond_Lattimore
Richmond Pearson Hobson	http://en.wikipedia.org/wiki/Richmond_Pearson_Hobson
Rick Allen	http://en.wikipedia.org/wiki/Rick_Allen_(drummer)
Rick Boucher	http://en.wikipedia.org/wiki/Rick_Boucher
Rick Boucher	http://en.wikipedia.org/wiki/Rick_Boucher
Rick Danko	http://en.wikipedia.org/wiki/Rick_Danko
Rick Dees	http://en.wikipedia.org/wiki/Rick_Dees
Rick Derringer	http://en.wikipedia.org/wiki/Rick_Derringer
Rick Fox	http://en.wikipedia.org/wiki/Rick_Fox
Rick Hall	http://en.wikipedia.org/wiki/Rick_Hall
Rick Hurst	http://en.wikipedia.org/wiki/Rick_Hurst
Rick James	http://en.wikipedia.org/wiki/Rick_James
Rick Jason	http://en.wikipedia.org/wiki/Rick_Jason
Rick Kemp	http://en.wikipedia.org/wiki/Rick_Kemp
Rick Larsen	http://en.wikipedia.org/wiki/Rick_Larsen
Rick Lazio	http://en.wikipedia.org/wiki/Rick_Lazio
Rick Majerus	http://en.wikipedia.org/wiki/Rick_Majerus
Rick Mears	http://en.wikipedia.org/wiki/Rick_Mears
Rick Metsger	http://en.wikipedia.org/wiki/Rick_Metsger
Rick Moody	http://en.wikipedia.org/wiki/Rick_Moody
Rick Moranis	http://en.wikipedia.org/wiki/Rick_Moranis
Rick Perry	http://en.wikipedia.org/wiki/Rick_Perry
Rick Perry	http://en.wikipedia.org/wiki/Rick_Perry
Rick Renzi	http://en.wikipedia.org/wiki/Rick_Renzi
Rick Rescorla	http://en.wikipedia.org/wiki/Rick_Rescorla
Rick Ross	http://en.wikipedia.org/wiki/Rick_Ross_(consultant)
Rick Rubin	http://en.wikipedia.org/wiki/Rick_Rubin
Rick Santorum	http://en.wikipedia.org/wiki/Rick_Santorum
Rick Savage	http://en.wikipedia.org/wiki/Rick_Savage
Rick Scarborough	http://en.wikipedia.org/wiki/Rick_Scarborough
Rick Schroder	http://en.wikipedia.org/wiki/Rick_Schroder
Rick Smith	http://en.wikipedia.org/wiki/Rick_Smith_%28American_football%29
Rick Springfield	http://en.wikipedia.org/wiki/Rick_Springfield
Rick Stephens	http://en.wikipedia.org/wiki/Rick_Stephens
Rick Wagoner	http://en.wikipedia.org/wiki/Rick_Wagoner
Rick Wakeman	http://en.wikipedia.org/wiki/Rick_Wakeman
Rick Warren	http://en.wikipedia.org/wiki/Rick_Warren
Rick Wright	http://en.wikipedia.org/wiki/Rick_Wright
Rickey Henderson	http://en.wikipedia.org/wiki/Rickey_Henderson
Ricki Lake	http://en.wikipedia.org/wiki/Ricki_Lake
Rickie Lee Jones	http://en.wikipedia.org/wiki/Rickie_Lee_Jones
Ricky Gervais	http://en.wikipedia.org/wiki/Ricky_Gervais
Ricky Martin	http://en.wikipedia.org/wiki/Ricky_Martin
Ricky Nelson	http://en.wikipedia.org/wiki/Ricky_Nelson
Ricky Ponting	http://en.wikipedia.org/wiki/Ricky_Ponting
Ricky Skaggs	http://en.wikipedia.org/wiki/Ricky_Skaggs
Ricky Ullman	http://en.wikipedia.org/wiki/Ricky_Ullman
Ricky Williams	http://en.wikipedia.org/wiki/Ricky_Williams
Ricky Wilson	http://en.wikipedia.org/wiki/Ricky_Wilson_(American_musician)
Rider Strong	http://en.wikipedia.org/wiki/Rider_Strong
Ridley Scott	http://en.wikipedia.org/wiki/Ridley_Scott
Rigoberta Mench� Tum	http://en.wikipedia.org/wiki/Rigoberta_Mench%FA_Tum
Rik Mayall	http://en.wikipedia.org/wiki/Rik_Mayall
Riki Rachtman	http://en.wikipedia.org/wiki/Riki_Rachtman
Rikki Fulton	http://en.wikipedia.org/wiki/Rikki_Fulton
Riley Smith	http://en.wikipedia.org/wiki/Riley_Smith
Ring Lardner	http://en.wikipedia.org/wiki/Ring_Lardner
Ring Lardner, Jr.	http://en.wikipedia.org/wiki/Ring_Lardner%2C_Jr.
Ringo Starr	http://en.wikipedia.org/wiki/Ringo_Starr
Rio Ferdinand	http://en.wikipedia.org/wiki/Rio_Ferdinand
Rip Taylor	http://en.wikipedia.org/wiki/Rip_Taylor
Rip Torn	http://en.wikipedia.org/wiki/Rip_Torn
Rita Coolidge	http://en.wikipedia.org/wiki/Rita_Coolidge
Rita Cosby	http://en.wikipedia.org/wiki/Rita_Cosby
Rita Dove	http://en.wikipedia.org/wiki/Rita_Dove
Rita Hayworth	http://en.wikipedia.org/wiki/Rita_Hayworth
Rita Mae Brown	http://en.wikipedia.org/wiki/Rita_Mae_Brown
Rita Moreno	http://en.wikipedia.org/wiki/Rita_Moreno
Rita Rudner	http://en.wikipedia.org/wiki/Rita_Rudner
Rita Wilson	http://en.wikipedia.org/wiki/Rita_Wilson
Ritchie Barrett	http://en.wikipedia.org/wiki/Richard_Barrett_(musician)
Ritchie Blackmore	http://en.wikipedia.org/wiki/Ritchie_Blackmore
Ritchie Valens	http://en.wikipedia.org/wiki/Ritchie_Valens
River Phoenix	http://en.wikipedia.org/wiki/River_Phoenix
Rivers Cuomo	http://en.wikipedia.org/wiki/Rivers_Cuomo
Rjyan Kidwell	http://en.wikipedia.org/wiki/Rjyan_Kidwell
Roald Amundsen	http://en.wikipedia.org/wiki/Roald_Amundsen
Roald Dahl	http://en.wikipedia.org/wiki/Roald_Dahl
Roald Hoffmann	http://en.wikipedia.org/wiki/Roald_Hoffmann
Rob "CmdrTaco" Malda	http://en.wikipedia.org/wiki/Rob_Malda
Rob Bishop	http://en.wikipedia.org/wiki/Rob_Bishop
Rob Bourdon	http://en.wikipedia.org/wiki/Rob_Bourdon
Rob Brown	http://en.wikipedia.org/wiki/Rob_Brown_(actor)
Rob Brown	http://en.wikipedia.org/wiki/Rob_Brown_(musician)
Rob Corddry	http://en.wikipedia.org/wiki/Rob_Corddry
Rob Dibble	http://en.wikipedia.org/wiki/Rob_Dibble
Rob Estes	http://en.wikipedia.org/wiki/Rob_Estes
Rob Glaser	http://en.wikipedia.org/wiki/Rob_Glaser
Rob Halford	http://en.wikipedia.org/wiki/Rob_Halford
Rob Liefeld	http://en.wikipedia.org/wiki/Rob_Liefeld
Rob Lowe	http://en.wikipedia.org/wiki/Rob_Lowe
Rob Morrow	http://en.wikipedia.org/wiki/Rob_Morrow
Rob Pilatus	http://en.wikipedia.org/wiki/Rob_Pilatus
Rob Portman	http://en.wikipedia.org/wiki/Rob_Portman
Rob Reiner	http://en.wikipedia.org/wiki/Rob_Reiner
Rob Schneider	http://en.wikipedia.org/wiki/Rob_Schneider
Rob Simmons	http://en.wikipedia.org/wiki/Rob_Simmons
Rob Thomas	http://en.wikipedia.org/wiki/Rob_Thomas_(musician)
Rob Walton	http://en.wikipedia.org/wiki/Rob_Walton
Rob Wexler	http://en.wikipedia.org/wiki/Rob_Wexler
Rob Wilson	http://en.wikipedia.org/wiki/Rob_Wilson
Rob Wittman	http://en.wikipedia.org/wiki/Rob_Wittman
Rob Zombie	http://en.wikipedia.org/wiki/Rob_Zombie
Robbie Coltrane	http://en.wikipedia.org/wiki/Robbie_Coltrane
Robbie Fowler	http://en.wikipedia.org/wiki/Robbie_Fowler
Robbie Knievel	http://en.wikipedia.org/wiki/Robbie_Knievel
Robbie Robertson	http://en.wikipedia.org/wiki/Robbie_Robertson
Robbie Williams	http://en.wikipedia.org/wiki/Robbie_Williams
Robby Benson	http://en.wikipedia.org/wiki/Robby_Benson
Robby Krieger	http://en.wikipedia.org/wiki/Robby_Krieger
Robert A. Borski	http://en.wikipedia.org/wiki/Robert_A._Borski
Robert A. Heinlein	http://en.wikipedia.org/wiki/Robert_A._Heinlein
Robert A. Lovett	http://en.wikipedia.org/wiki/Robert_A._Lovett
Robert A. Millikan	http://en.wikipedia.org/wiki/Robert_A._Millikan
Robert A. Mundell	http://en.wikipedia.org/wiki/Robert_A._Mundell
Robert A. Roe	http://en.wikipedia.org/wiki/Robert_A._Roe
Robert A. Taft	http://en.wikipedia.org/wiki/Robert_A._Taft
Robert A. Young	http://en.wikipedia.org/wiki/Robert_A._Young
Robert Adam	http://en.wikipedia.org/wiki/Robert_Adam
Robert Aderholt	http://en.wikipedia.org/wiki/Robert_Aderholt
Robert Alda	http://en.wikipedia.org/wiki/Robert_Alda
Robert Aldrich	http://en.wikipedia.org/wiki/Robert_Aldrich
Robert Allston	http://en.wikipedia.org/wiki/Robert_Allston
Robert Altman	http://en.wikipedia.org/wiki/Robert_Altman
Robert Ambrose	http://en.wikipedia.org/wiki/Robert_Ambrose_%28conductor%29
Robert Anton Wilson	http://en.wikipedia.org/wiki/Robert_Anton_Wilson
Robert Arthur Talbot Gascoyne-Cecil	http://en.wikipedia.org/wiki/Robert_Arthur_Talbot_Gascoyne-Cecil
Robert Asprin	http://en.wikipedia.org/wiki/Robert_Asprin
Robert Atkins	http://en.wikipedia.org/wiki/Robert_Atkins_(nutritionist)
Robert B. Laughlin	http://en.wikipedia.org/wiki/Robert_B._Laughlin
Robert B. Silvers	http://en.wikipedia.org/wiki/Robert_B._Silvers
Robert B. Woodward	http://en.wikipedia.org/wiki/Robert_B._Woodward
Robert Bacon	http://en.wikipedia.org/wiki/Robert_Bacon
Robert Baden-Powell	http://en.wikipedia.org/wiki/Robert_Baden-Powell
Robert Baer	http://en.wikipedia.org/wiki/Robert_Baer
Robert Bakewell	http://en.wikipedia.org/wiki/Robert_Bakewell_(agriculturalist)
Robert Barnes	http://en.wikipedia.org/wiki/Robert_Barnes_(martyr)
Robert Bellarmine	http://en.wikipedia.org/wiki/Robert_Bellarmine
Robert Beltran	http://en.wikipedia.org/wiki/Robert_Beltran
Robert Benchley	http://en.wikipedia.org/wiki/Robert_Benchley
Robert Bennett	http://en.wikipedia.org/wiki/Bob_Bennett_(politician)
Robert Benton	http://en.wikipedia.org/wiki/Robert_Benton
Robert Blake	http://en.wikipedia.org/wiki/Robert_Blake_(actor)
Robert Bly	http://en.wikipedia.org/wiki/Robert_Bly
Robert Bolt	http://en.wikipedia.org/wiki/Robert_Bolt
Robert Bork	http://en.wikipedia.org/wiki/Robert_Bork
Robert Boyle	http://en.wikipedia.org/wiki/Robert_Boyle
Robert Brady	http://en.wikipedia.org/wiki/Bob_Brady
Robert Bresson	http://en.wikipedia.org/wiki/Robert_Bresson
Robert Bridges	http://en.wikipedia.org/wiki/Robert_Bridges
Robert Brown	http://en.wikipedia.org/wiki/Robert_Brown_(botanist)
Robert Browning	http://en.wikipedia.org/wiki/Robert_Browning
Robert Brustein	http://en.wikipedia.org/wiki/Robert_Brustein
Robert Buckland	http://en.wikipedia.org/wiki/Robert_Buckland
Robert Burns	http://en.wikipedia.org/wiki/Robert_Burns
Robert Burton	http://en.wikipedia.org/wiki/Robert_Burton_(scholar)
Robert Byrd	http://en.wikipedia.org/wiki/Robert_Byrd
Robert C. Byrd	http://en.wikipedia.org/wiki/Robert_C._Byrd
Robert C. Gallo	http://en.wikipedia.org/wiki/Robert_C._Gallo
Robert C. Merton	http://en.wikipedia.org/wiki/Robert_C._Merton
Robert C. Richardson	http://en.wikipedia.org/wiki/Robert_Coleman_Richardson
Robert C. Smith	http://en.wikipedia.org/wiki/Robert_C._Smith
Robert Cantwell	http://en.wikipedia.org/wiki/Robert_Cantwell
Robert Carlyle	http://en.wikipedia.org/wiki/Robert_Carlyle
Robert Caro	http://en.wikipedia.org/wiki/Robert_Caro
Robert Carradine	http://en.wikipedia.org/wiki/Robert_Carradine
Robert Cecil	http://en.wikipedia.org/wiki/Robert_Cecil,_1st_Viscount_Cecil_of_Chelwood
Robert Chambers	http://en.wikipedia.org/wiki/Robert_Chambers
Robert Charles Winthrop	http://en.wikipedia.org/wiki/Robert_Charles_Winthrop
Robert Clary	http://en.wikipedia.org/wiki/Robert_Clary
Robert Clive	http://en.wikipedia.org/wiki/Robert_Clive
Robert Conrad	http://en.wikipedia.org/wiki/Robert_Conrad
Robert Cormier	http://en.wikipedia.org/wiki/Robert_Cormier
Robert Cotton	http://en.wikipedia.org/wiki/Robert_Bruce_Cotton
Robert Cray	http://en.wikipedia.org/wiki/Robert_Cray
Robert Creeley	http://en.wikipedia.org/wiki/Robert_Creeley
Robert Crippen	http://en.wikipedia.org/wiki/Robert_Crippen
Robert Crumb	http://en.wikipedia.org/wiki/Robert_Crumb
Robert Culp	http://en.wikipedia.org/wiki/Robert_Culp
Robert Cutler	http://en.wikipedia.org/wiki/Robert_Cutler
Robert D. Kaplan	http://en.wikipedia.org/wiki/Robert_D._Kaplan
Robert D. McEwen	http://en.wikipedia.org/wiki/Robert_D._McEwen
Robert D. Steele	http://en.wikipedia.org/wiki/Robert_D._Steele
Robert D. Walter	http://en.wikipedia.org/wiki/Robert_D._Walter
Robert Dale Owen	http://en.wikipedia.org/wiki/Robert_Dale_Owen
Robert De Niro	http://en.wikipedia.org/wiki/Robert_De_Niro
Robert del Naja	http://en.wikipedia.org/wiki/Robert_del_Naja
Robert Donat	http://en.wikipedia.org/wiki/Robert_Donat
Robert Downey, Jr.	http://en.wikipedia.org/wiki/Robert_Downey%2C_Jr.
Robert Downey, Sr.	http://en.wikipedia.org/wiki/Robert_Downey%2C_Sr.
Robert Drinan	http://en.wikipedia.org/wiki/Robert_Drinan
Robert Duncan	http://en.wikipedia.org/wiki/Robert_Duncan_(poet)
Robert Duvall	http://en.wikipedia.org/wiki/Robert_Duvall
Robert E. Andrews	http://en.wikipedia.org/wiki/Robert_E._Andrews
Robert E. Badham	http://en.wikipedia.org/wiki/Robert_E._Badham
Robert E. Howard	http://en.wikipedia.org/wiki/Robert_E._Howard
Robert E. Kahn	http://en.wikipedia.org/wiki/Robert_E._Kahn
Robert E. Lee	http://en.wikipedia.org/wiki/Robert_E._Lee
Robert E. Park	http://en.wikipedia.org/wiki/Robert_E._Park
Robert E. Peary	http://en.wikipedia.org/wiki/Robert_E._Peary
Robert E. Rubin	http://en.wikipedia.org/wiki/Robert_E._Rubin
Robert E. Sherwood	http://en.wikipedia.org/wiki/Robert_E._Sherwood
Robert E. Smylie	http://en.wikipedia.org/wiki/Robert_E._Smylie
Robert E. Wise, Jr.	http://en.wikipedia.org/wiki/Robert_E._Wise%2C_Jr.
Robert Ehrlich	http://en.wikipedia.org/wiki/Robert_Ehrlich
Robert Englund	http://en.wikipedia.org/wiki/Robert_Englund
Robert Evans	http://en.wikipedia.org/wiki/Robert_Evans_(producer)
Robert F. Curl, Jr.	http://en.wikipedia.org/wiki/Robert_F._Curl%2C_Jr.
Robert F. Ellsworth	http://en.wikipedia.org/wiki/Robert_F._Ellsworth
Robert F. Kennedy	http://en.wikipedia.org/wiki/Robert_F._Kennedy
Robert F. Kennedy, Jr.	http://en.wikipedia.org/wiki/Robert_F._Kennedy%2C_Jr.
Robert F. Smith	http://en.wikipedia.org/wiki/Robert_F._Smith
Robert F. Wagner, Jr.	http://en.wikipedia.org/wiki/Robert_F._Wagner%2C_Jr.
Robert F. Wagner, Sr.	http://en.wikipedia.org/wiki/Robert_F._Wagner
Robert Fico	http://en.wikipedia.org/wiki/Robert_Fico
Robert Fisk	http://en.wikipedia.org/wiki/Robert_Fisk
Robert Flello	http://en.wikipedia.org/wiki/Robert_Flello
Robert Fludd	http://en.wikipedia.org/wiki/Robert_Fludd
Robert Forster	http://en.wikipedia.org/wiki/Robert_Forster
Robert Foxworth	http://en.wikipedia.org/wiki/Robert_Foxworth
Robert Fripp	http://en.wikipedia.org/wiki/Robert_Fripp
Robert Frost	http://en.wikipedia.org/wiki/Robert_Frost
Robert Fuller	http://en.wikipedia.org/wiki/Robert_Fuller_(actor)
Robert Fuller	http://en.wikipedia.org/wiki/Robert_Fuller
Robert Fulton	http://en.wikipedia.org/wiki/Robert_Fulton
Robert G. Ingersoll	http://en.wikipedia.org/wiki/Robert_G._Ingersoll
Robert G. Torricelli	http://en.wikipedia.org/wiki/Robert_G._Torricelli
Robert Gant	http://en.wikipedia.org/wiki/Robert_Gant
Robert Garcia	http://en.wikipedia.org/wiki/Robert_García
Robert Garioch	http://en.wikipedia.org/wiki/Robert_Garioch
Robert Garnier	http://en.wikipedia.org/wiki/Robert_Garnier
Robert Gates	http://en.wikipedia.org/wiki/Robert_Gates
Robert Giaimo	http://en.wikipedia.org/wiki/Robert_Giaimo
Robert Gibbs	http://en.wikipedia.org/wiki/Robert_Gibbs
Robert Goddard	http://en.wikipedia.org/wiki/Robert_Goddard
Robert Goodwill	http://en.wikipedia.org/wiki/Robert_Goodwill
Robert Goulet	http://en.wikipedia.org/wiki/Robert_Goulet
Robert Grant	http://en.wikipedia.org/wiki/Robert_Grant_(novelist)
Robert Graves	http://en.wikipedia.org/wiki/Robert_Graves
Robert Greene	http://en.wikipedia.org/wiki/Robert_Greene_(dramatist)
Robert Greenwald	http://en.wikipedia.org/wiki/Robert_Greenwald
Robert Greifeld	http://en.wikipedia.org/wiki/Robert_Greifeld
Robert Grosseteste	http://en.wikipedia.org/wiki/Robert_Grosseteste
Robert Guillaume	http://en.wikipedia.org/wiki/Robert_Guillaume
Robert Guiscard	http://en.wikipedia.org/wiki/Robert_Guiscard
Robert H. Jackson	http://en.wikipedia.org/wiki/Robert_H._Jackson
Robert H. Michel	http://en.wikipedia.org/wiki/Robert_H._Michel
Robert Halfon	http://en.wikipedia.org/wiki/Robert_Halfon
Robert Hamerling	http://en.wikipedia.org/wiki/Robert_Hamerling
Robert Hanssen	http://en.wikipedia.org/wiki/Robert_Hanssen
Robert Hass	http://en.wikipedia.org/wiki/Robert_Hass
Robert Hawke	http://en.wikipedia.org/wiki/Robert_Hawke
Robert Hayden	http://en.wikipedia.org/wiki/Robert_Hayden
Robert Hays	http://en.wikipedia.org/wiki/Robert_Hays
Robert Heilbroner	http://en.wikipedia.org/wiki/Robert_Heilbroner
Robert Herrick	http://en.wikipedia.org/wiki/Robert_Herrick_(poet)
Robert Hill	http://en.wikipedia.org/wiki/Robert_Hill_(Australian_diplomat)
Robert Hofstadter	http://en.wikipedia.org/wiki/Robert_Hofstadter
Robert Hooke	http://en.wikipedia.org/wiki/Robert_Hooke
Robert Hossein	http://en.wikipedia.org/wiki/Robert_Hossein
Robert Huber	http://en.wikipedia.org/wiki/Robert_Huber
Robert I	http://en.wikipedia.org/wiki/Robert_I_of_France
Robert Iger	http://en.wikipedia.org/wiki/Robert_Iger
Robert II	http://en.wikipedia.org/wiki/Robert_II_of_France
Robert III	http://en.wikipedia.org/wiki/Robert_III
Robert Iler	http://en.wikipedia.org/wiki/Robert_Iler
Robert Indiana	http://en.wikipedia.org/wiki/Robert_Indiana
Robert J. Aumann	http://en.wikipedia.org/wiki/Robert_J._Aumann
Robert J. Lagomarsino	http://en.wikipedia.org/wiki/Robert_J._Lagomarsino
Robert J. Mrazek	http://en.wikipedia.org/wiki/Robert_J._Mrazek
Robert Jarvik	http://en.wikipedia.org/wiki/Robert_Jarvik
Robert Jenkins	http://en.wikipedia.org/wiki/Robert_Jenkins_(master_mariner)
Robert Johnson	http://en.wikipedia.org/wiki/Robert_Johnson_(musician)
Robert Jordan	http://en.wikipedia.org/wiki/Robert_Jordan
Robert K. Dornan	http://en.wikipedia.org/wiki/Robert_K._Dornan
Robert K. Merton	http://en.wikipedia.org/wiki/Robert_K._Merton
Robert K. Ressler	http://en.wikipedia.org/wiki/Robert_K._Ressler
Robert Kagan	http://en.wikipedia.org/wiki/Robert_Kagan
Robert Kardashian	http://en.wikipedia.org/wiki/Robert_Kardashian
Robert Keable	http://en.wikipedia.org/wiki/Robert_Keable
Robert Kiyosaki	http://en.wikipedia.org/wiki/Robert_Kiyosaki
Robert Klein	http://en.wikipedia.org/wiki/Robert_Klein
Robert Koch	http://en.wikipedia.org/wiki/Robert_Koch
Robert Kocharyan	http://en.wikipedia.org/wiki/Robert_Kocharyan
Robert Kraft	http://en.wikipedia.org/wiki/Robert_Kraft
Robert L. Johnson	http://en.wikipedia.org/wiki/Robert_L._Johnson
Robert L. Livingston Jr.	http://en.wikipedia.org/wiki/Bob_Livingston
Robert L. Ripley	http://en.wikipedia.org/wiki/Robert_L._Ripley
Robert Laird Borden	http://en.wikipedia.org/wiki/Robert_Laird_Borden
Robert Lansing	http://en.wikipedia.org/wiki/Robert_Lansing
Robert Latham Owen	http://en.wikipedia.org/wiki/Robert_Latham_Owen
Robert Leighton	http://en.wikipedia.org/wiki/Robert_Leighton_(prelate)
Robert Lewis Taylor	http://en.wikipedia.org/wiki/Robert_Lewis_Taylor
Robert Ley	http://en.wikipedia.org/wiki/Robert_Ley
Robert Lindsay	http://en.wikipedia.org/wiki/Robert_Lindsay_(actor)
Robert List	http://en.wikipedia.org/wiki/Robert_List
Robert Loggia	http://en.wikipedia.org/wiki/Robert_Loggia
Robert Louis Stevenson	http://en.wikipedia.org/wiki/Robert_Louis_Stevenson
Robert Lowell	http://en.wikipedia.org/wiki/Robert_Lowell
Robert Lowery	http://en.wikipedia.org/wiki/Robert_Lowery_(actor)
Robert Lucas	http://en.wikipedia.org/wiki/Robert_Lucas,_Jr.
Robert Ludlum	http://en.wikipedia.org/wiki/Robert_Ludlum
Robert Luskin	http://en.wikipedia.org/wiki/Robert_Luskin
Robert M. Gates	http://en.wikipedia.org/wiki/Robert_M._Gates
Robert M. Solow	http://en.wikipedia.org/wiki/Robert_M._Solow
Robert MacNeil	http://en.wikipedia.org/wiki/Robert_MacNeil
Robert Mannyng	http://en.wikipedia.org/wiki/Robert_Mannyng
Robert Mapplethorpe	http://en.wikipedia.org/wiki/Robert_Mapplethorpe
Robert Mathews	http://en.wikipedia.org/wiki/Robert_Jay_Mathews
Robert Matsui	http://en.wikipedia.org/wiki/Robert_Matsui
Robert McAlmon	http://en.wikipedia.org/wiki/Robert_McAlmon
Robert McNamara	http://en.wikipedia.org/wiki/Robert_McNamara
Robert Menendez	http://en.wikipedia.org/wiki/Robert_Menendez
Robert Menzies	http://en.wikipedia.org/wiki/Robert_Menzies
Robert Mitchum	http://en.wikipedia.org/wiki/Robert_Mitchum
Robert Mondavi	http://en.wikipedia.org/wiki/Robert_Mondavi
Robert Montgomery	http://en.wikipedia.org/wiki/Robert_Montgomery_(actor)
Robert Moog	http://en.wikipedia.org/wiki/Robert_Moog
Robert Morley	http://en.wikipedia.org/wiki/Robert_Morley
Robert Morris	http://en.wikipedia.org/wiki/Robert_Morris_(financier)
Robert Morris, Jr.	http://en.wikipedia.org/wiki/Robert_Tappan_Morris
Robert Morrison MacIver	http://en.wikipedia.org/wiki/Robert_Morrison_MacIver
Robert Morse	http://en.wikipedia.org/wiki/Robert_Morse
Robert Mosbacher	http://en.wikipedia.org/wiki/Robert_Mosbacher
Robert Moses	http://en.wikipedia.org/wiki/Robert_Moses
Robert Mueller	http://en.wikipedia.org/wiki/Robert_Mueller
Robert Mugabe	http://en.wikipedia.org/wiki/Robert_Mugabe
Robert Mulligan	http://en.wikipedia.org/wiki/Robert_Mulligan
Robert Musil	http://en.wikipedia.org/wiki/Robert_Musil
Robert Newton	http://en.wikipedia.org/wiki/Robert_Newton
Robert Noel	http://en.wikipedia.org/wiki/Robert_Noel
Robert Novak	http://en.wikipedia.org/wiki/Robert_Novak
Robert Nozick	http://en.wikipedia.org/wiki/Robert_Nozick
Robert O. Bowen	http://en.wikipedia.org/wiki/Robert_O._Bowen
Robert of Clermont	http://en.wikipedia.org/wiki/Robert,_Count_of_Clermont
Robert O'Hara Burke	http://en.wikipedia.org/wiki/Robert_O%27Hara_Burke
Robert Olen Butler	http://en.wikipedia.org/wiki/Robert_Olen_Butler
Robert Oppenheimer	http://en.wikipedia.org/wiki/Robert_Oppenheimer
Robert Orben	http://en.wikipedia.org/wiki/Robert_Orben
Robert Owen	http://en.wikipedia.org/wiki/Robert_Owen
Robert P. Casey	http://en.wikipedia.org/wiki/Robert_P._Casey
Robert P. Tristram Coffin	http://en.wikipedia.org/wiki/Robert_P._Tristram_Coffin
Robert Palmer	http://en.wikipedia.org/wiki/Robert_Palmer_(singer)
Robert Papp	http://en.wikipedia.org/wiki/Robert_Papp
Robert Parish	http://en.wikipedia.org/wiki/Robert_Parish
Robert Pastorelli	http://en.wikipedia.org/wiki/Robert_Pastorelli
Robert Patrick	http://en.wikipedia.org/wiki/Robert_Patrick
Robert Peel	http://en.wikipedia.org/wiki/Robert_Peel
Robert Penn Warren	http://en.wikipedia.org/wiki/Robert_Penn_Warren
Robert Picardo	http://en.wikipedia.org/wiki/Robert_Picardo
Robert Pickton	http://en.wikipedia.org/wiki/Robert_Pickton
Robert Pinsky	http://en.wikipedia.org/wiki/Robert_Pinsky
Robert Plant	http://en.wikipedia.org/wiki/Robert_Plant
Robert Powell	http://en.wikipedia.org/wiki/Robert_Powell
Robert Preston	http://en.wikipedia.org/wiki/Robert_Preston_(actor)
Robert Quine	http://en.wikipedia.org/wiki/Robert_Quine
Robert R. Livingston	http://en.wikipedia.org/wiki/Robert_Livingston_(1746–1813)
Robert Rauschenberg	http://en.wikipedia.org/wiki/Robert_Rauschenberg
Robert Redford	http://en.wikipedia.org/wiki/Robert_Redford
Robert Reed	http://en.wikipedia.org/wiki/Robert_Reed
Robert Reich	http://en.wikipedia.org/wiki/Robert_Reich
Robert Riley	http://en.wikipedia.org/wiki/Bob_C._Riley
Robert Rodriguez	http://en.wikipedia.org/wiki/Robert_Rodriguez
Robert Runcie	http://en.wikipedia.org/wiki/Robert_Runcie
Robert Ryan	http://en.wikipedia.org/wiki/Robert_Ryan
Robert S. Brookings	http://en.wikipedia.org/wiki/Robert_S._Brookings
Robert S. Mulliken	http://en.wikipedia.org/wiki/Robert_S._Mulliken
Robert S. Strauss	http://en.wikipedia.org/wiki/Robert_S._Strauss
Robert Scheer	http://en.wikipedia.org/wiki/Robert_Scheer
Robert Schrieffer	http://en.wikipedia.org/wiki/Robert_Schrieffer
Robert Schuller	http://en.wikipedia.org/wiki/Robert_Schuller
Robert Schumann	http://en.wikipedia.org/wiki/Robert_Schumann
Robert Sean Leonard	http://en.wikipedia.org/wiki/Robert_Sean_Leonard
Robert Shapiro	http://en.wikipedia.org/wiki/Robert_Shapiro_(lawyer)
Robert Shaw	http://en.wikipedia.org/wiki/Robert_Shaw_(actor)
Robert Shaye	http://en.wikipedia.org/wiki/Robert_Shaye
Robert Shea	http://en.wikipedia.org/wiki/Robert_Shea
Robert Silverberg	http://en.wikipedia.org/wiki/Robert_Silverberg
Robert Smigel	http://en.wikipedia.org/wiki/Robert_Smigel
Robert Smith	http://en.wikipedia.org/wiki/Sir_Robert_Smith,_3rd_Baronet
Robert Smith	http://en.wikipedia.org/wiki/Robert_Smith_(musician)
Robert Smith Surtees	http://en.wikipedia.org/wiki/Robert_Smith_Surtees
Robert Smith Walker	http://en.wikipedia.org/wiki/Robert_Smith_Walker
Robert Southey	http://en.wikipedia.org/wiki/Robert_Southey
Robert Stack	http://en.wikipedia.org/wiki/Robert_Stack
Robert Stephenson	http://en.wikipedia.org/wiki/Robert_Stephenson
Robert Sterling	http://en.wikipedia.org/wiki/Robert_Sterling
Robert Stevenson	http://en.wikipedia.org/wiki/Robert_Stevenson_(civil_engineer)
Robert Stevenson	http://en.wikipedia.org/wiki/Robert_Stevenson_(director)
Robert Stewart, Viscount Castlereagh	http://en.wikipedia.org/wiki/Robert_Stewart%2C_Viscount_Castlereagh
Robert Stone	http://en.wikipedia.org/wiki/Robert_Stone_(novelist)
Robert Surtees	http://en.wikipedia.org/wiki/Robert_Surtees_(antiquarian)
Robert Syms	http://en.wikipedia.org/wiki/Robert_Syms
Robert T. Bakker	http://en.wikipedia.org/wiki/Robert_T._Bakker
Robert T. Matsui	http://en.wikipedia.org/wiki/Robert_T._Matsui
Robert T. Stafford	http://en.wikipedia.org/wiki/Robert_T._Stafford
Robert Taylor	http://en.wikipedia.org/wiki/Robert_Taylor_(actor)
Robert the Bruce	http://en.wikipedia.org/wiki/Robert_the_Bruce
Robert Thorne	http://en.wikipedia.org/wiki/Robert_Thorne
Robert Tilton	http://en.wikipedia.org/wiki/Robert_Tilton
Robert Todd Lincoln	http://en.wikipedia.org/wiki/Robert_Todd_Lincoln
Robert Torricelli	http://en.wikipedia.org/wiki/Robert_Torricelli
Robert Towne	http://en.wikipedia.org/wiki/Robert_Towne
Robert Townsend	http://en.wikipedia.org/wiki/Robert_Townsend_(actor)
Robert Trimble	http://en.wikipedia.org/wiki/Robert_Trimble
Robert Trujillo	http://en.wikipedia.org/wiki/Robert_Trujillo
Robert Urich	http://en.wikipedia.org/wiki/Robert_Urich
Robert Vaughn	http://en.wikipedia.org/wiki/Robert_Vaughn
Robert Venturi	http://en.wikipedia.org/wiki/Robert_Venturi
Robert W. Anderson	http://en.wikipedia.org/wiki/Robert_W._Anderson
Robert W. Davis	http://en.wikipedia.org/wiki/Robert_William_Davis
Robert W. Kastenmeier	http://en.wikipedia.org/wiki/Robert_W._Kastenmeier
Robert W. Service	http://en.wikipedia.org/wiki/Robert_W._Service
Robert W. Tucker	http://en.wikipedia.org/wiki/Robert_W._Tucker
Robert W. Wood	http://en.wikipedia.org/wiki/Robert_W._Wood
Robert Wagner	http://en.wikipedia.org/wiki/Robert_Wagner
Robert Walker	http://en.wikipedia.org/wiki/Robert_Walker_(actor)
Robert Walpole	http://en.wikipedia.org/wiki/Robert_Walpole
Robert Walter	http://en.wikipedia.org/wiki/Robert_Walter
Robert Wilhelm Bunsen	http://en.wikipedia.org/wiki/Robert_Wilhelm_Bunsen
Robert Wilson	http://en.wikipedia.org/wiki/Robert_Wilson_(director)
Robert Wise	http://en.wikipedia.org/wiki/Robert_Wise
Robert Woodrow Wilson	http://en.wikipedia.org/wiki/Robert_Woodrow_Wilson
Robert Wuhl	http://en.wikipedia.org/wiki/Robert_Wuhl
Robert Wyatt	http://en.wikipedia.org/wiki/Robert_Wyatt
Robert X. Cringely	http://en.wikipedia.org/wiki/Robert_X._Cringely
Robert Young	http://en.wikipedia.org/wiki/Robert_Young_(actor)
Robert Z. Leonard	http://en.wikipedia.org/wiki/Robert_Z._Leonard
Robert Zemeckis	http://en.wikipedia.org/wiki/Robert_Zemeckis
Roberta Blackman-Woods	http://en.wikipedia.org/wiki/Roberta_Blackman-Woods
Roberta Flack	http://en.wikipedia.org/wiki/Roberta_Flack
Roberta Williams	http://en.wikipedia.org/wiki/Roberta_Williams
Robert-Fran�ois Damiens	http://en.wikipedia.org/wiki/Robert-Fran%E7ois_Damiens
Roberto Alomar	http://en.wikipedia.org/wiki/Roberto_Alomar
Roberto Baggio	http://en.wikipedia.org/wiki/Roberto_Baggio
Roberto Benigni	http://en.wikipedia.org/wiki/Roberto_Benigni
Roberto Calvi	http://en.wikipedia.org/wiki/Roberto_Calvi
Roberto Carlos	http://en.wikipedia.org/wiki/Roberto_Carlos_(singer)
Roberto Cavalli	http://en.wikipedia.org/wiki/Roberto_Cavalli
Roberto Clemente	http://en.wikipedia.org/wiki/Roberto_Clemente
Roberto Duran	http://en.wikipedia.org/wiki/Roberto_Duran
Roberto Mangabeira Unger	http://en.wikipedia.org/wiki/Roberto_Mangabeira_Unger
Roberto Rossellini	http://en.wikipedia.org/wiki/Roberto_Rossellini
Robertson Davies	http://en.wikipedia.org/wiki/Robertson_Davies
Robin Cook	http://en.wikipedia.org/wiki/Robin_Cook_(American_novelist)
Robin Cook	http://en.wikipedia.org/wiki/Robin_Cook
Robin Gibb	http://en.wikipedia.org/wiki/Robin_Gibb
Robin Givens	http://en.wikipedia.org/wiki/Robin_Givens
Robin Guthrie	http://en.wikipedia.org/wiki/Robin_Guthrie
Robin Hayes	http://en.wikipedia.org/wiki/Robin_Hayes
Robin Leach	http://en.wikipedia.org/wiki/Robin_Leach
Robin McKinley	http://en.wikipedia.org/wiki/Robin_McKinley
Robin Quivers	http://en.wikipedia.org/wiki/Robin_Quivers
Robin Roberts	http://en.wikipedia.org/wiki/Robin_Roberts_(newscaster)
Robin Roberts	http://en.wikipedia.org/wiki/Robin_Roberts_(baseball)
Robin Tallon	http://en.wikipedia.org/wiki/Robin_Tallon
Robin Trower	http://en.wikipedia.org/wiki/Robin_Trower
Robin Tunney	http://en.wikipedia.org/wiki/Robin_Tunney
Robin Walker	http://en.wikipedia.org/wiki/Robin_Walker_(politician)
Robin Williams	http://en.wikipedia.org/wiki/Robin_Williams
Robin Wright Penn	http://en.wikipedia.org/wiki/Robin_Wright_Penn
Robin Yount	http://en.wikipedia.org/wiki/Robin_Yount
Robin Zander	http://en.wikipedia.org/wiki/Robin_Zander
Robinson Jeffers	http://en.wikipedia.org/wiki/Robinson_Jeffers
Robyn Hitchcock	http://en.wikipedia.org/wiki/Robyn_Hitchcock
Rocco DiSpirito	http://en.wikipedia.org/wiki/Rocco_DiSpirito
Rock Hudson	http://en.wikipedia.org/wiki/Rock_Hudson
Rockwell Kent	http://en.wikipedia.org/wiki/Rockwell_Kent
Rocky Graziano	http://en.wikipedia.org/wiki/Rocky_Graziano
Rocky Marciano	http://en.wikipedia.org/wiki/Rocky_Marciano
Rod Argent	http://en.wikipedia.org/wiki/Rod_Argent
Rod Blagojevich	http://en.wikipedia.org/wiki/Rod_Blagojevich
Rod Blagojevich	http://en.wikipedia.org/wiki/Rod_Blagojevich
Rod Carew	http://en.wikipedia.org/wiki/Rod_Carew
Rod Chandler	http://en.wikipedia.org/wiki/Rod_Chandler
Rod Chandler	http://en.wikipedia.org/wiki/Rod_Chandler
Rod Laver	http://en.wikipedia.org/wiki/Rod_Laver
Rod McKuen	http://en.wikipedia.org/wiki/Rod_McKuen
Rod Paige	http://en.wikipedia.org/wiki/Rod_Paige
Rod Serling	http://en.wikipedia.org/wiki/Rod_Serling
Rod Steiger	http://en.wikipedia.org/wiki/Rod_Steiger
Rod Stewart	http://en.wikipedia.org/wiki/Rod_Stewart
Rod Taylor	http://en.wikipedia.org/wiki/Rod_Taylor
Rodd Keith	http://en.wikipedia.org/wiki/Rodd_Keith
Roddy Doyle	http://en.wikipedia.org/wiki/Roddy_Doyle
Roddy McDowall	http://en.wikipedia.org/wiki/Roddy_McDowall
Roddy Piper	http://en.wikipedia.org/wiki/Roddy_Piper
Roderick MacKinnon	http://en.wikipedia.org/wiki/Roderick_MacKinnon
Rodney Alexander	http://en.wikipedia.org/wiki/Rodney_Alexander
Rodney Allen Rippy	http://en.wikipedia.org/wiki/Rodney_Allen_Rippy
Rodney Dangerfield	http://en.wikipedia.org/wiki/Rodney_Dangerfield
Rodney Frelinghuysen	http://en.wikipedia.org/wiki/Rodney_Frelinghuysen
Rodney King	http://en.wikipedia.org/wiki/Rodney_King
Rodney Slater	http://en.wikipedia.org/wiki/Rodney_E._Slater
Rodolphe T�pffer	http://en.wikipedia.org/wiki/Rodolphe_T%F6pffer
Rodrigo Rato	http://en.wikipedia.org/wiki/Rodrigo_Rato
Rodrigo Santoro	http://en.wikipedia.org/wiki/Rodrigo_Santoro
Roger Abbott	http://en.wikipedia.org/wiki/Roger_Abbott
Roger Adams	http://en.wikipedia.org/wiki/Roger_Adams
Roger Ailes	http://en.wikipedia.org/wiki/Roger_Ailes
Roger Alborough	http://en.wikipedia.org/wiki/Roger_Alborough
Roger Allam	http://en.wikipedia.org/wiki/Roger_Allam
Roger Ascham	http://en.wikipedia.org/wiki/Roger_Ascham
Roger Avary	http://en.wikipedia.org/wiki/Roger_Avary
Roger Babson	http://en.wikipedia.org/wiki/Roger_Babson
Roger Bacon	http://en.wikipedia.org/wiki/Roger_Bacon
Roger Bannister	http://en.wikipedia.org/wiki/Roger_Bannister
Roger Bart	http://en.wikipedia.org/wiki/Roger_Bart
Roger Boyle	http://en.wikipedia.org/wiki/Roger_Boyle
Roger Brooke Taney	http://en.wikipedia.org/wiki/Roger_Brooke_Taney
Roger Casement	http://en.wikipedia.org/wiki/Roger_Casement
Roger Clemens	http://en.wikipedia.org/wiki/Roger_Clemens
Roger Clinton	http://en.wikipedia.org/wiki/Roger_Clinton,_Jr.
Roger Cook	http://en.wikipedia.org/wiki/Roger_Cook_(landscaper)
Roger Corman	http://en.wikipedia.org/wiki/Roger_Corman
Roger Craig	http://en.wikipedia.org/wiki/Roger_Craig_(American_football)
Roger Daltrey	http://en.wikipedia.org/wiki/Roger_Daltrey
Roger E. Mosley	http://en.wikipedia.org/wiki/Roger_E._Mosley
Roger Ebert	http://en.wikipedia.org/wiki/Roger_Ebert
Roger Federer	http://en.wikipedia.org/wiki/Roger_Federer
Roger Gale	http://en.wikipedia.org/wiki/Roger_Gale
Roger Godsiff	http://en.wikipedia.org/wiki/Roger_Godsiff
Roger Hargreaves	http://en.wikipedia.org/wiki/Roger_Hargreaves
Roger Lodge	http://en.wikipedia.org/wiki/Roger_Lodge
Roger Mahony	http://en.wikipedia.org/wiki/Roger_Mahony
Roger Maris	http://en.wikipedia.org/wiki/Roger_Maris
Roger McGuinn	http://en.wikipedia.org/wiki/Roger_McGuinn
Roger Miller	http://en.wikipedia.org/wiki/Roger_Miller
Roger Moore	http://en.wikipedia.org/wiki/Roger_Moore
Roger Mudd	http://en.wikipedia.org/wiki/Roger_Mudd
Roger Nordlund	http://en.wikipedia.org/wiki/Roger_Nordlund
Roger Penrose	http://en.wikipedia.org/wiki/Roger_Penrose
Roger Sant	http://en.wikipedia.org/wiki/Roger_Sant
Roger Sessions	http://en.wikipedia.org/wiki/Roger_Sessions
Roger Sherman	http://en.wikipedia.org/wiki/Roger_Sherman
Roger Smith	http://en.wikipedia.org/wiki/Roger_Smith_(executive)
Roger Spottiswoode	http://en.wikipedia.org/wiki/Roger_Spottiswoode
Roger Staubach	http://en.wikipedia.org/wiki/Roger_Staubach
Roger Stone	http://en.wikipedia.org/wiki/Roger_Stone
Roger Taylor	http://en.wikipedia.org/wiki/Roger_Taylor_(Duran_Duran_drummer)
Roger Taylor	http://en.wikipedia.org/wiki/Roger_Meddows-Taylor
Roger Tubby	http://en.wikipedia.org/wiki/Roger_Tubby
Roger Vadim	http://en.wikipedia.org/wiki/Roger_Vadim
Roger Waters	http://en.wikipedia.org/wiki/Roger_Waters
Roger Wicker	http://en.wikipedia.org/wiki/Roger_Wicker
Roger Wilkins	http://en.wikipedia.org/wiki/Roger_Wilkins
Roger Williams	http://en.wikipedia.org/wiki/Roger_Williams_(UK_politician)
Roger Williams	http://en.wikipedia.org/wiki/Roger_Williams_(theologian)
Roger Zelazny	http://en.wikipedia.org/wiki/Roger_Zelazny
Rogers C.B. Morton	http://en.wikipedia.org/wiki/Rogers_C.B._Morton
Rogers Hornsby	http://en.wikipedia.org/wiki/Rogers_Hornsby
Rogier van der Weyden	http://en.wikipedia.org/wiki/Rogier_van_der_Weyden
Roh Moo Hyun	http://en.wikipedia.org/wiki/Roh_Moo_Hyun
Roh Moo-hyun	http://en.wikipedia.org/wiki/Roh_Moo-hyun
Roh Tae Woo	http://en.wikipedia.org/wiki/Roh_Tae_Woo
Rokusaburo Michiba	http://en.wikipedia.org/wiki/Rokusaburo_Michiba
Roky Erickson	http://en.wikipedia.org/wiki/Roky_Erickson
Roland Barthes	http://en.wikipedia.org/wiki/Roland_Barthes
Roland Burris	http://en.wikipedia.org/wiki/Roland_Burris
Roland Culver	http://en.wikipedia.org/wiki/Roland_Culver
Roland Emmerich	http://en.wikipedia.org/wiki/Roland_Emmerich
Roland Freisler	http://en.wikipedia.org/wiki/Roland_Freisler
Roland Gift	http://en.wikipedia.org/wiki/Roland_Gift
Roland Joff�	http://en.wikipedia.org/wiki/Roland_Joff%E9
Roland Martin	http://en.wikipedia.org/wiki/Roland_Martin_(fisherman)
Rollen Stewart	http://en.wikipedia.org/wiki/Rollen_Stewart
Rollie Fingers	http://en.wikipedia.org/wiki/Rollie_Fingers
Rollo May	http://en.wikipedia.org/wiki/Rollo_May
Roma Downey	http://en.wikipedia.org/wiki/Roma_Downey
Roma Maffia	http://en.wikipedia.org/wiki/Roma_Maffia
Romain Rolland	http://en.wikipedia.org/wiki/Romain_Rolland
Roman Cieslewicz	http://en.wikipedia.org/wiki/Roman_Cieslewicz
Roman Gabriel	http://en.wikipedia.org/wiki/Roman_Gabriel
Roman Herzog	http://en.wikipedia.org/wiki/Roman_Herzog
Roman Hruska	http://en.wikipedia.org/wiki/Roman_Hruska
Roman Polanski	http://en.wikipedia.org/wiki/Roman_Polanski
Romano L. Mazzoli	http://en.wikipedia.org/wiki/Romano_L._Mazzoli
Romano Prodi	http://en.wikipedia.org/wiki/Romano_Prodi
Romano Prodi	http://en.wikipedia.org/wiki/Romano_Prodi
Romare Bearden	http://en.wikipedia.org/wiki/Romare_Bearden
Romolo Valli	http://en.wikipedia.org/wiki/Romolo_Valli
Romy Schneider	http://en.wikipedia.org/wiki/Romy_Schneider
Ron Artest	http://en.wikipedia.org/wiki/Ron_Artest
Ron Atkinson	http://en.wikipedia.org/wiki/Ron_Atkinson
Ron Brown	http://en.wikipedia.org/wiki/Ron_Brown_(U.S._politician)
Ron Burkle	http://en.wikipedia.org/wiki/Ron_Burkle
Ron Burton	http://en.wikipedia.org/wiki/Ron_Burton
Ron Carey	http://en.wikipedia.org/wiki/Ron_Carey_(labor_leader)
Ron Chernow	http://en.wikipedia.org/wiki/Ron_Chernow
Ron Davies	http://en.wikipedia.org/wiki/Ron_Davies_%28Welsh_politician%29
Ron de Lugo	http://en.wikipedia.org/wiki/Ron_de_Lugo
Ron Dellums	http://en.wikipedia.org/wiki/Ron_Dellums
Ron Eldard	http://en.wikipedia.org/wiki/Ron_Eldard
Ron Ely	http://en.wikipedia.org/wiki/Ron_Ely
Ron Geesin	http://en.wikipedia.org/wiki/Ron_Geesin
Ron Glass	http://en.wikipedia.org/wiki/Ron_Glass
Ron Howard	http://en.wikipedia.org/wiki/Ron_Howard
Ron Kind	http://en.wikipedia.org/wiki/Ron_Kind
Ron Klein	http://en.wikipedia.org/wiki/Ron_Klein
Ron Klink	http://en.wikipedia.org/wiki/Ron_Klink
Ron Leibman	http://en.wikipedia.org/wiki/Ron_Leibman
Ron Lewis	http://en.wikipedia.org/wiki/Ron_Lewis
Ron Livingston	http://en.wikipedia.org/wiki/Ron_Livingston
Ron Marlenee	http://en.wikipedia.org/wiki/Ron_Marlenee
Ron McKernan	http://en.wikipedia.org/wiki/Ron_McKernan
Ron Moody	http://en.wikipedia.org/wiki/Ron_Moody
Ron Nessen	http://en.wikipedia.org/wiki/Ron_Nessen
Ron O'Neal	http://en.wikipedia.org/wiki/Ron_O%27Neal
Ron Packard	http://en.wikipedia.org/wiki/Ron_Packard
Ron Palillo	http://en.wikipedia.org/wiki/Ron_Palillo
Ron Paul	http://en.wikipedia.org/wiki/Ron_Paul
Ron Perelman	http://en.wikipedia.org/wiki/Ron_Perelman
Ron Perlman	http://en.wikipedia.org/wiki/Ron_Perlman
Ron Popeil	http://en.wikipedia.org/wiki/Ron_Popeil
Ron Reagan	http://en.wikipedia.org/wiki/Ron_Reagan
Ron Santo	http://en.wikipedia.org/wiki/Ron_Santo
Ron Silver	http://en.wikipedia.org/wiki/Ron_Silver
Ron Suskind	http://en.wikipedia.org/wiki/Ron_Suskind
Ron Weaver	http://en.wikipedia.org/wiki/Ron_Weaver
Ron White	http://en.wikipedia.org/wiki/Ron_White
Ron Wood	http://en.wikipedia.org/wiki/Ron_Wood
Ron Wyden	http://en.wikipedia.org/wiki/Ron_Wyden
Ron Wyden	http://en.wikipedia.org/wiki/Ron_Wyden
Ron Ziegler	http://en.wikipedia.org/wiki/Ron_Ziegler
Rona Barrett	http://en.wikipedia.org/wiki/Rona_Barrett
Rona Jaffe	http://en.wikipedia.org/wiki/Rona_Jaffe
Ronald Cohen	http://en.wikipedia.org/wiki/Ronald_Cohen
Ronald Colman	http://en.wikipedia.org/wiki/Ronald_Colman
Ronald D. Coleman	http://en.wikipedia.org/wiki/Ronald_D._Coleman
Ronald D. Sugar	http://en.wikipedia.org/wiki/Ronald_Sugar
Ronald Dworkin	http://en.wikipedia.org/wiki/Ronald_Dworkin
Ronald G. W. Norrish	http://en.wikipedia.org/wiki/Ronald_G._W._Norrish
Ronald H. Coase	http://en.wikipedia.org/wiki/Ronald_H._Coase
Ronald Isley	http://en.wikipedia.org/wiki/Ronald_Isley
Ronald Neame	http://en.wikipedia.org/wiki/Ronald_Neame
Ronald Reagan	http://en.wikipedia.org/wiki/Ronald_Reagan
Ronald Ross	http://en.wikipedia.org/wiki/Ronald_Ross
Ronald Steel	http://en.wikipedia.org/wiki/Ronald_Steel
Ronald V. Dellums	http://en.wikipedia.org/wiki/Ronald_V._Dellums
Ronald Venetiaan	http://en.wikipedia.org/wiki/Ronald_Venetiaan
Ronaldinho	http://en.wikipedia.org/wiki/Ronaldinho
Ronan Keating	http://en.wikipedia.org/wiki/Ronan_Keating
Roni Size	http://en.wikipedia.org/wiki/Roni_Size
Ronn Moss	http://en.wikipedia.org/wiki/Ronn_Moss
Ronn Owens	http://en.wikipedia.org/wiki/Ronn_Owens
Ronnie Barker	http://en.wikipedia.org/wiki/Ronnie_Barker
Ronnie Biggs	http://en.wikipedia.org/wiki/Ronnie_Biggs
Ronnie Campbell	http://en.wikipedia.org/wiki/Ronnie_Campbell
Ronnie Corbett	http://en.wikipedia.org/wiki/Ronnie_Corbett
Ronnie Earle	http://en.wikipedia.org/wiki/Ronnie_Earle
Ronnie G. Flippo	http://en.wikipedia.org/wiki/Ronnie_G._Flippo
Ronnie James Dio	http://en.wikipedia.org/wiki/Ronnie_James_Dio
Ronnie Milsap	http://en.wikipedia.org/wiki/Ronnie_Milsap
Ronnie Montrose	http://en.wikipedia.org/wiki/Ronnie_Montrose
Ronnie Musgrove	http://en.wikipedia.org/wiki/Ronnie_Musgrove
Ronnie Spector	http://en.wikipedia.org/wiki/Ronnie_Spector
Ronnie Van Zant	http://en.wikipedia.org/wiki/Ronnie_Van_Zant
Ronnie White	http://en.wikipedia.org/wiki/Ronnie_White
Ronny Cox	http://en.wikipedia.org/wiki/Ronny_Cox
Roone Arledge	http://en.wikipedia.org/wiki/Roone_Arledge
Roosevelt Skerrit	http://en.wikipedia.org/wiki/Roosevelt_Skerrit
Roots Manuva	http://en.wikipedia.org/wiki/Roots_Manuva
Rory Calhoun	http://en.wikipedia.org/wiki/Rory_Calhoun
Rory Cochrane	http://en.wikipedia.org/wiki/Rory_Cochrane
Rory Culkin	http://en.wikipedia.org/wiki/Rory_Culkin
Rory Stewart	http://en.wikipedia.org/wiki/Rory_Stewart
Rosa Blasi	http://en.wikipedia.org/wiki/Rosa_Blasi
Rosa DeLauro	http://en.wikipedia.org/wiki/Rosa_DeLauro
Rosa Luxemburg	http://en.wikipedia.org/wiki/Rosa_Luxemburg
Rosa Parks	http://en.wikipedia.org/wiki/Rosa_Parks
Rosalind Cash	http://en.wikipedia.org/wiki/Rosalind_Cash
Rosalind Chao	http://en.wikipedia.org/wiki/Rosalind_Chao
Rosalind Russell	http://en.wikipedia.org/wiki/Rosalind_Russell
Rosalyn Sussman Yalow	http://en.wikipedia.org/wiki/Rosalyn_Sussman_Yalow
Rosalynn Carter	http://en.wikipedia.org/wiki/Rosalynn_Carter
Rosamund Pike	http://en.wikipedia.org/wiki/Rosamund_Pike
Rosanna Arquette	http://en.wikipedia.org/wiki/Rosanna_Arquette
Rosanne Cash	http://en.wikipedia.org/wiki/Rosanne_Cash
Rosario Dawson	http://en.wikipedia.org/wiki/Rosario_Dawson
Roscoe Bartlett	http://en.wikipedia.org/wiki/Roscoe_Bartlett
Roscoe Conkling	http://en.wikipedia.org/wiki/Roscoe_Conkling
Roscoe H. Hillenkoetter	http://en.wikipedia.org/wiki/Roscoe_H._Hillenkoetter
Roscoe Mitchell	http://en.wikipedia.org/wiki/Roscoe_Mitchell
Roscoe Pound	http://en.wikipedia.org/wiki/Roscoe_Pound
Rose Abdoo	http://en.wikipedia.org/wiki/Rose_Abdoo
Rose Hobart	http://en.wikipedia.org/wiki/Rose_Hobart
Rose Kennedy	http://en.wikipedia.org/wiki/Rose_Kennedy
Rose Marie	http://en.wikipedia.org/wiki/Rose_Marie
Rose Mary Woods	http://en.wikipedia.org/wiki/Rose_Mary_Woods
Rose McGowan	http://en.wikipedia.org/wiki/Rose_McGowan
Roseanne Barr	http://en.wikipedia.org/wiki/Roseanne_Barr
Roselyn Sanchez	http://en.wikipedia.org/wiki/Roselyn_Sanchez
Rosemary Clooney	http://en.wikipedia.org/wiki/Rosemary_Clooney
Rosemary Harris	http://en.wikipedia.org/wiki/Rosemary_Harris
Rosemary Kennedy	http://en.wikipedia.org/wiki/Rosemary_Kennedy
Rosemary Murphy	http://en.wikipedia.org/wiki/Rosemary_Murphy
Rosemary West	http://en.wikipedia.org/wiki/Rosemary_West
Rosey Grier	http://en.wikipedia.org/wiki/Rosey_Grier
Roshumba Williams	http://en.wikipedia.org/wiki/Roshumba_Williams
Rosie Cooper	http://en.wikipedia.org/wiki/Rosie_Cooper
Rosie O'Donnell	http://en.wikipedia.org/wiki/Rosie_O%27Donnell
Rosie Perez	http://en.wikipedia.org/wiki/Rosie_Perez
Rosie Winterton	http://en.wikipedia.org/wiki/Rosie_Winterton
Ross Alexander	http://en.wikipedia.org/wiki/Ross_Alexander
Ross Bagdasarian	http://en.wikipedia.org/wiki/Ross_Bagdasarian,_Sr.
Ross Macdonald	http://en.wikipedia.org/wiki/Ross_Macdonald
Ross Martin	http://en.wikipedia.org/wiki/Ross_Martin
Ross McElwee	http://en.wikipedia.org/wiki/Ross_McElwee
Ross McWhirter	http://en.wikipedia.org/wiki/Ross_McWhirter
Rossano Brazzi	http://en.wikipedia.org/wiki/Rossano_Brazzi
Rouben Mamoulian	http://en.wikipedia.org/wiki/Rouben_Mamoulian
Rowan Atkinson	http://en.wikipedia.org/wiki/Rowan_Atkinson
Rowan Scarborough	http://en.wikipedia.org/wiki/Rowan_Scarborough
Rowan Williams	http://en.wikipedia.org/wiki/Rowan_Williams
Rowland Evans	http://en.wikipedia.org/wiki/Rowland_Evans
Roxanne Hart	http://en.wikipedia.org/wiki/Roxanne_Hart
Roxanne Shante	http://en.wikipedia.org/wiki/Roxanne_Shante
Roxie Roker	http://en.wikipedia.org/wiki/Roxie_Roker
Roy Acuff	http://en.wikipedia.org/wiki/Roy_Acuff
Roy Barnes	http://en.wikipedia.org/wiki/Roy_Barnes
Roy Blount, Jr.	http://en.wikipedia.org/wiki/Roy_Blount%2C_Jr.
Roy Blunt	http://en.wikipedia.org/wiki/Roy_Blunt
Roy Campanella	http://en.wikipedia.org/wiki/Roy_Campanella
Roy Clark	http://en.wikipedia.org/wiki/Roy_Clark
Roy Cohn	http://en.wikipedia.org/wiki/Roy_Cohn
Roy D. Chapin, Jr.	http://en.wikipedia.org/wiki/Roy_D._Chapin%2C_Jr.
Roy D. Chapin, Sr.	http://en.wikipedia.org/wiki/Roy_D._Chapin
Roy Del Ruth	http://en.wikipedia.org/wiki/Roy_Del_Ruth
Roy Dyson	http://en.wikipedia.org/wiki/Roy_Dyson
Roy E. Disney	http://en.wikipedia.org/wiki/Roy_E._Disney
Roy Eldridge	http://en.wikipedia.org/wiki/Roy_Eldridge
Roy Harper	http://en.wikipedia.org/wiki/Roy_Harper
Roy Harrod	http://en.wikipedia.org/wiki/Roy_Harrod
Roy Horn	http://en.wikipedia.org/wiki/Roy_Horn
Roy Hudd	http://en.wikipedia.org/wiki/Roy_Hudd
Roy Innis	http://en.wikipedia.org/wiki/Roy_Innis
Roy Keane	http://en.wikipedia.org/wiki/Roy_Keane
Roy Lee Johnson	http://en.wikipedia.org/wiki/Roy_Lee_Johnson
Roy Lichtenstein	http://en.wikipedia.org/wiki/Roy_Lichtenstein
Roy Moore	http://en.wikipedia.org/wiki/Roy_Moore
Roy O. Disney	http://en.wikipedia.org/wiki/Roy_O._Disney
Roy Orbison	http://en.wikipedia.org/wiki/Roy_Orbison
Roy Rogers	http://en.wikipedia.org/wiki/Roy_Rogers
Roy Romer	http://en.wikipedia.org/wiki/Roy_Romer
Roy Scheider	http://en.wikipedia.org/wiki/Roy_Scheider
Roy Welensky	http://en.wikipedia.org/wiki/Roy_Welensky
Roy William Neill	http://en.wikipedia.org/wiki/Roy_William_Neill
Roy Williams	http://en.wikipedia.org/wiki/Roy_Williams_(artist)
Roy Wood	http://en.wikipedia.org/wiki/Roy_Wood
Royal Rife	http://en.wikipedia.org/wiki/Royal_Rife
Royall Tyler	http://en.wikipedia.org/wiki/Royall_Tyler
Roza Otunbayeva	http://en.wikipedia.org/wiki/Roza_Otunbayeva
Rozanne L. Ridgway	http://en.wikipedia.org/wiki/Rozanne_L._Ridgway
Rozonda "Chilli" Thomas	http://en.wikipedia.org/wiki/Rozonda_%22Chilli%22_Thomas
Rube Goldberg	http://en.wikipedia.org/wiki/Rube_Goldberg
Ruben Blades	http://en.wikipedia.org/wiki/Ruben_Blades
Rub�n Dar�o	http://en.wikipedia.org/wiki/Rub%E9n_Dar%EDo
Rub�n Hinojosa	http://en.wikipedia.org/wiki/Rub%E9n_Hinojosa
Ruben Salazar	http://en.wikipedia.org/wiki/Ruben_Salazar
Ruben Studdard	http://en.wikipedia.org/wiki/Ruben_Studdard
Ruby Dee	http://en.wikipedia.org/wiki/Ruby_Dee
Ruby Keeler	http://en.wikipedia.org/wiki/Ruby_Keeler
Rudolf Carnap	http://en.wikipedia.org/wiki/Rudolf_Carnap
Rudolf Clausius	http://en.wikipedia.org/wiki/Rudolf_Clausius
Rudolf Diesel	http://en.wikipedia.org/wiki/Rudolf_Diesel
Rudolf Eucken	http://en.wikipedia.org/wiki/Rudolf_Eucken
Rudolf Hess	http://en.wikipedia.org/wiki/Rudolf_Hess
Rudolf M�ssbauer	http://en.wikipedia.org/wiki/Rudolf_M%F6ssbauer
Rudolf Nureyev	http://en.wikipedia.org/wiki/Rudolf_Nureyev
Rudolf Peierls	http://en.wikipedia.org/wiki/Rudolf_Peierls
Rudolf Schenker	http://en.wikipedia.org/wiki/Rudolf_Schenker
Rudolf Schuster	http://en.wikipedia.org/wiki/Rudolf_Schuster
Rudolfo Anaya	http://en.wikipedia.org/wiki/Rudolfo_Anaya
Rudolph A. Marcus	http://en.wikipedia.org/wiki/Rudolph_A._Marcus
Rudolph Valentino	http://en.wikipedia.org/wiki/Rudolph_Valentino
Rudy Bond	http://en.wikipedia.org/wiki/Rudy_Bond
Rudy Boschwitz	http://en.wikipedia.org/wiki/Rudy_Boschwitz
Rudy Giuliani	http://en.wikipedia.org/wiki/Rudy_Giuliani
Rudy Rucker	http://en.wikipedia.org/wiki/Rudy_Rucker
Rudy Tomjanovich	http://en.wikipedia.org/wiki/Rudy_Tomjanovich
Rudy Vallee	http://en.wikipedia.org/wiki/Rudy_Vallee
Rudyard Kipling	http://en.wikipedia.org/wiki/Rudyard_Kipling
Rue McClanahan	http://en.wikipedia.org/wiki/Rue_McClanahan
Rufino Tamayo	http://en.wikipedia.org/wiki/Rufino_Tamayo
Rufus Choate	http://en.wikipedia.org/wiki/Rufus_Choate
Rufus Putnam	http://en.wikipedia.org/wiki/Rufus_Putnam
Rufus Sewell	http://en.wikipedia.org/wiki/Rufus_Sewell
Rufus Wainwright	http://en.wikipedia.org/wiki/Rufus_Wainwright
Ruggero Giuseppe Boscovich	http://en.wikipedia.org/wiki/Ruggero_Giuseppe_Boscovich
Ruggero Leoncavallo	http://en.wikipedia.org/wiki/Ruggero_Leoncavallo
Rula Lenska	http://en.wikipedia.org/wiki/Rula_Lenska
Rupert Brooke	http://en.wikipedia.org/wiki/Rupert_Brooke
Rupert Everett	http://en.wikipedia.org/wiki/Rupert_Everett
Rupert Graves	http://en.wikipedia.org/wiki/Rupert_Graves
Rupert Grint	http://en.wikipedia.org/wiki/Rupert_Grint
Rupert Holmes	http://en.wikipedia.org/wiki/Rupert_Holmes
Rupert Murdoch	http://en.wikipedia.org/wiki/Rupert_Murdoch
Rupert Sheldrake	http://en.wikipedia.org/wiki/Rupert_Sheldrake
Rupiah Banda	http://en.wikipedia.org/wiki/Rupiah_Banda
Rush Holt	http://en.wikipedia.org/wiki/Rush_Holt
Rush Limbaugh	http://en.wikipedia.org/wiki/Rush_Limbaugh
Rushanara Ali	http://en.wikipedia.org/wiki/Rushanara_Ali
Rushdy Abaza	http://en.wikipedia.org/wiki/Rushdy_Abaza
Russ Abbot	http://en.wikipedia.org/wiki/Russ_Abbot
Russ Carnahan	http://en.wikipedia.org/wiki/Russ_Carnahan
Russ Feingold	http://en.wikipedia.org/wiki/Russ_Feingold
Russ Meyer	http://en.wikipedia.org/wiki/Russ_Meyer
Russ Morgan	http://en.wikipedia.org/wiki/Russ_Morgan
Russ Tamblyn	http://en.wikipedia.org/wiki/Russ_Tamblyn
Russel Crouse	http://en.wikipedia.org/wiki/Russel_Crouse
Russel Honore	http://en.wikipedia.org/wiki/Russel_Honore
Russell A. Alger	http://en.wikipedia.org/wiki/Russell_A._Alger
Russell A. Hulse	http://en.wikipedia.org/wiki/Russell_A._Hulse
Russell B. Long	http://en.wikipedia.org/wiki/Russell_B._Long
Russell Baker	http://en.wikipedia.org/wiki/Russell_Baker
Russell Banks	http://en.wikipedia.org/wiki/Russell_Banks
Russell Boyd	http://en.wikipedia.org/wiki/Russell_Boyd
Russell Brown	http://en.wikipedia.org/wiki/Russell_Brown
Russell Crowe	http://en.wikipedia.org/wiki/Russell_Crowe
Russell Hitchcock	http://en.wikipedia.org/wiki/Russell_Hitchcock
Russell Hunter	http://en.wikipedia.org/wiki/Russell_Hunter
Russell Johnson	http://en.wikipedia.org/wiki/Russell_Johnson
Russell Johnson	http://en.wikipedia.org/wiki/Russell_Johnson
Russell Kirk	http://en.wikipedia.org/wiki/Russell_Kirk
Russell Simmons	http://en.wikipedia.org/wiki/Russell_Simmons
Russell Simmons	http://en.wikipedia.org/wiki/Russell_Simmons
Russell W. Peterson	http://en.wikipedia.org/wiki/Russell_W._Peterson
Russell Wong	http://en.wikipedia.org/wiki/Russell_Wong
Rusty Cundieff	http://en.wikipedia.org/wiki/Rusty_Cundieff
Rusty Schweickart	http://en.wikipedia.org/wiki/Rusty_Schweickart
Rutger Hauer	http://en.wikipedia.org/wiki/Rutger_Hauer
Ruth Ann Minner	http://en.wikipedia.org/wiki/Ruth_Ann_Minner
Ruth Ann Minner	http://en.wikipedia.org/wiki/Ruth_Ann_Minner
Ruth Bader Ginsburg	http://en.wikipedia.org/wiki/Ruth_Bader_Ginsburg
Ruth Benedict	http://en.wikipedia.org/wiki/Ruth_Benedict
Ruth Brown	http://en.wikipedia.org/wiki/Ruth_Brown
Ruth Bryan Owen	http://en.wikipedia.org/wiki/Ruth_Bryan_Owen
Ruth Buzzi	http://en.wikipedia.org/wiki/Ruth_Buzzi
Ruth Chatterton	http://en.wikipedia.org/wiki/Ruth_Chatterton
Ruth Ellis	http://en.wikipedia.org/wiki/Ruth_Ellis
Ruth Ford	http://en.wikipedia.org/wiki/Ruth_Ford_(actress)
Ruth Gordon	http://en.wikipedia.org/wiki/Ruth_Gordon
Ruth Hussey	http://en.wikipedia.org/wiki/Ruth_Hussey
Ruth Lilly	http://en.wikipedia.org/wiki/Ruth_Lilly
Ruth McDevitt	http://en.wikipedia.org/wiki/Ruth_McDevitt
Ruth McKenney	http://en.wikipedia.org/wiki/Ruth_McKenney
Ruth Parasol	http://en.wikipedia.org/wiki/Ruth_Parasol
Ruth Pointer	http://en.wikipedia.org/wiki/Ruth_Pointer
Ruth Porter Crawford	http://en.wikipedia.org/wiki/Ruth_Porter_Crawford
Ruth Prawer Jhabvala	http://en.wikipedia.org/wiki/Ruth_Prawer_Jhabvala
Ruth Underwood	http://en.wikipedia.org/wiki/Ruth_Underwood
Ruth Warrick	http://en.wikipedia.org/wiki/Ruth_Warrick
Ruth Westheimer	http://en.wikipedia.org/wiki/Ruth_Westheimer
Rutherford B. Hayes	http://en.wikipedia.org/wiki/Rutherford_B._Hayes
Ruud Gullit	http://en.wikipedia.org/wiki/Ruud_Gullit
Ruud van Nistelrooy	http://en.wikipedia.org/wiki/Ruud_van_Nistelrooy
Ruy Teixeira	http://en.wikipedia.org/wiki/Ruy_Teixeira
Ry Cooder	http://en.wikipedia.org/wiki/Ry_Cooder
Ryan Adams	http://en.wikipedia.org/wiki/Ryan_Adams
Ryan Cabrera	http://en.wikipedia.org/wiki/Ryan_Cabrera
Ryan Carnes	http://en.wikipedia.org/wiki/Ryan_Carnes
Ryan Dunn	http://en.wikipedia.org/wiki/Ryan_Dunn
Ryan Giggs	http://en.wikipedia.org/wiki/Ryan_Giggs
Ryan Gosling	http://en.wikipedia.org/wiki/Ryan_Gosling
Ryan Merriman	http://en.wikipedia.org/wiki/Ryan_Merriman
Ryan Murphy	http://en.wikipedia.org/wiki/Ryan_Murphy_(writer)
Ryan O'Neal	http://en.wikipedia.org/wiki/Ryan_O%27Neal
Ryan Phillippe	http://en.wikipedia.org/wiki/Ryan_Phillippe
Ryan Reynolds	http://en.wikipedia.org/wiki/Ryan_Reynolds
Ryan Seacrest	http://en.wikipedia.org/wiki/Ryan_Seacrest
Ryan Stiles	http://en.wikipedia.org/wiki/Ryan_Stiles
Ryan White	http://en.wikipedia.org/wiki/Ryan_White
Ryoji Noyori	http://en.wikipedia.org/wiki/Ryoji_Noyori
Ryszard Kuklinski	http://en.wikipedia.org/wiki/Ryszard_Kuklinski
Ryutaro Hashimoto	http://en.wikipedia.org/wiki/Ryutaro_Hashimoto
S. E. Hinton	http://en.wikipedia.org/wiki/S._E._Hinton
S. Epatha Merkerson	http://en.wikipedia.org/wiki/S._Epatha_Merkerson
S. I. Hayakawa	http://en.wikipedia.org/wiki/S._I._Hayakawa
S. J. Perelman	http://en.wikipedia.org/wiki/S._J._Perelman
S. R. Nathan	http://en.wikipedia.org/wiki/S._R._Nathan
S. R. Nathan	http://en.wikipedia.org/wiki/S._R._Nathan
S. S. Van Dine	http://en.wikipedia.org/wiki/S._S._Van_Dine
S. Truett Cathy	http://en.wikipedia.org/wiki/S._Truett_Cathy
S. Weir Mitchell	http://en.wikipedia.org/wiki/S._Weir_Mitchell
S. William Green	http://en.wikipedia.org/wiki/S._William_Green
S.P. Somtow	http://en.wikipedia.org/wiki/S.P._Somtow
Saad Al-Abdullah Al-Salim Al-Sabah	http://en.wikipedia.org/wiki/Saad_Al-Abdullah_Al-Salim_Al-Sabah
Saad Hariri	http://en.wikipedia.org/wiki/Saad_Hariri
Sabah al-Ahmad al-Jabir al-Sabah	http://en.wikipedia.org/wiki/Sabah_al-Ahmad_al-Jabir_al-Sabah
Sabah IV al-Sabah	http://en.wikipedia.org/wiki/Sabah_Al-Ahmad_Al-Jaber_Al-Sabah
Sabrina LeBeauf	http://en.wikipedia.org/wiki/Sabrina_LeBeauf
Sabrina Lloyd	http://en.wikipedia.org/wiki/Sabrina_Lloyd
Sachin Tendulkar	http://en.wikipedia.org/wiki/Sachin_Tendulkar
Sadaharu Oh	http://en.wikipedia.org/wiki/Sadaharu_Oh
Saddam Hussein	http://en.wikipedia.org/wiki/Saddam_Hussein
Sadeq Hedayat	http://en.wikipedia.org/wiki/Sadeq_Hedayat
Sadi Carnot	http://en.wikipedia.org/wiki/Nicolas_Léonard_Sadi_Carnot
Sadie Frost	http://en.wikipedia.org/wiki/Sadie_Frost
Sadiq Khan	http://en.wikipedia.org/wiki/Sadiq_Khan
Saffron Burrows	http://en.wikipedia.org/wiki/Saffron_Burrows
Sai Baba	http://en.wikipedia.org/wiki/Sathya_Sai_Baba
Said Musa	http://en.wikipedia.org/wiki/Said_Musa
Saif al-Adel	http://en.wikipedia.org/wiki/Saif_al-Adel
Sait Faik Abasiyanik	http://en.wikipedia.org/wiki/Sait_Faik_Abasiyanik
Sajid Javid	http://en.wikipedia.org/wiki/Sajid_Javid
Sal Amendola	http://en.wikipedia.org/wiki/Sal_Amendola
Sal Mineo	http://en.wikipedia.org/wiki/Sal_Mineo
Sala Burton	http://en.wikipedia.org/wiki/Sala_Burton
Salem bin Laden	http://en.wikipedia.org/wiki/Salem_bin_Laden
Sali Berisha	http://en.wikipedia.org/wiki/Sali_Berisha
Sally Ann Howes	http://en.wikipedia.org/wiki/Sally_Ann_Howes
Sally Eastall	http://en.wikipedia.org/wiki/Sally_Eastall
Sally Eilers	http://en.wikipedia.org/wiki/Sally_Eilers
Sally Field	http://en.wikipedia.org/wiki/Sally_Field
Sally Hemings	http://en.wikipedia.org/wiki/Sally_Hemings
Sally Jessy Raphael	http://en.wikipedia.org/wiki/Sally_Jessy_Raphael
Sally Kellerman	http://en.wikipedia.org/wiki/Sally_Kellerman
Sally Kirkland	http://en.wikipedia.org/wiki/Sally_Kirkland
Sally Ride	http://en.wikipedia.org/wiki/Sally_Ride
Sally Struthers	http://en.wikipedia.org/wiki/Sally_Struthers
Salma Hayek	http://en.wikipedia.org/wiki/Salma_Hayek
Salman Khan	http://en.wikipedia.org/wiki/Salman_Khan
Salman Rushdie	http://en.wikipedia.org/wiki/Salman_Rushdie
Salmon P. Chase	http://en.wikipedia.org/wiki/Salmon_P._Chase
Salome Jens	http://en.wikipedia.org/wiki/Salome_Jens
Salou Djibo	http://en.wikipedia.org/wiki/Salou_Djibo
Salvador Allende	http://en.wikipedia.org/wiki/Salvador_Allende
Salvador Dali	http://en.wikipedia.org/wiki/Salvador_Dali
Salvador de Madariaga	http://en.wikipedia.org/wiki/Salvador_de_Madariaga
Salvador Luria	http://en.wikipedia.org/wiki/Salvador_Luria
Salvatore Maranzano	http://en.wikipedia.org/wiki/Salvatore_Maranzano
Salvatore Quasimodo	http://en.wikipedia.org/wiki/Salvatore_Quasimodo
Sam Beam	http://en.wikipedia.org/wiki/Sam_Beam
Sam Brown	http://en.wikipedia.org/wiki/Sam_Brown_(artist)
Sam Brownback	http://en.wikipedia.org/wiki/Sam_Brownback
Sam Champion	http://en.wikipedia.org/wiki/Sam_Champion
Sam Cooke	http://en.wikipedia.org/wiki/Sam_Cooke
Sam Dash	http://en.wikipedia.org/wiki/Sam_Dash
Sam Donaldson	http://en.wikipedia.org/wiki/Sam_Donaldson
Sam Elliott	http://en.wikipedia.org/wiki/Sam_Elliott
Sam Ervin	http://en.wikipedia.org/wiki/Sam_Ervin
Sam Farr	http://en.wikipedia.org/wiki/Sam_Farr
Sam Gejdenson	http://en.wikipedia.org/wiki/Sam_Gejdenson
Sam Giancana	http://en.wikipedia.org/wiki/Sam_Giancana
Sam Goddard	http://en.wikipedia.org/wiki/Sam_Goddard
Sam Graves	http://en.wikipedia.org/wiki/Sam_Graves
Sam Gyimah	http://en.wikipedia.org/wiki/Sam_Gyimah
Sam Hamm	http://en.wikipedia.org/wiki/Sam_Hamm
Sam Henderson	http://en.wikipedia.org/wiki/Sam_Henderson
Sam Hinds	http://en.wikipedia.org/wiki/Sam_Hinds
Sam Houston	http://en.wikipedia.org/wiki/Sam_Houston
Sam J. Jones	http://en.wikipedia.org/wiki/Sam_J._Jones
Sam Jaffe	http://en.wikipedia.org/wiki/Sam_Jaffe_(actor)
Sam Johnson	http://en.wikipedia.org/wiki/Sam_Johnson
Sam Kinison	http://en.wikipedia.org/wiki/Sam_Kinison
Sam M. Gibbons	http://en.wikipedia.org/wiki/Sam_M._Gibbons
Sam Mendes	http://en.wikipedia.org/wiki/Sam_Mendes
Sam Neill	http://en.wikipedia.org/wiki/Sam_Neill
Sam Nunn	http://en.wikipedia.org/wiki/Sam_Nunn
Sam Nunn	http://en.wikipedia.org/wiki/Sam_Nunn
Sam Palmisano	http://en.wikipedia.org/wiki/Sam_Palmisano
Sam Peckinpah	http://en.wikipedia.org/wiki/Sam_Peckinpah
Sam Phillips	http://en.wikipedia.org/wiki/Sam_Phillips
Sam Raimi	http://en.wikipedia.org/wiki/Sam_Raimi
Sam Rayburn	http://en.wikipedia.org/wiki/Sam_Rayburn
Sam Robards	http://en.wikipedia.org/wiki/Sam_Robards
Sam Rockwell	http://en.wikipedia.org/wiki/Sam_Rockwell
Sam Seder	http://en.wikipedia.org/wiki/Sam_Seder
Sam Shepard	http://en.wikipedia.org/wiki/Sam_Shepard
Sam Snead	http://en.wikipedia.org/wiki/Sam_Snead
Sam Tanenhaus	http://en.wikipedia.org/wiki/Sam_Tanenhaus
Sam Waksal	http://en.wikipedia.org/wiki/Sam_Waksal
Sam Walton	http://en.wikipedia.org/wiki/Sam_Walton
Sam Wanamaker	http://en.wikipedia.org/wiki/Sam_Wanamaker
Sam Waterston	http://en.wikipedia.org/wiki/Sam_Waterston
Sam Wood	http://en.wikipedia.org/wiki/Sam_Wood
Samaire Armstrong	http://en.wikipedia.org/wiki/Samaire_Armstrong
Samantha Bee	http://en.wikipedia.org/wiki/Samantha_Bee
Samantha Eggar	http://en.wikipedia.org/wiki/Samantha_Eggar
Samantha Mathis	http://en.wikipedia.org/wiki/Samantha_Mathis
Samantha Morton	http://en.wikipedia.org/wiki/Samantha_Morton
Samantha Mumba	http://en.wikipedia.org/wiki/Samantha_Mumba
Samantha Power	http://en.wikipedia.org/wiki/Samantha_Power
Samir Rifai	http://en.wikipedia.org/wiki/Samir_Rifai
Sammo Hung	http://en.wikipedia.org/wiki/Sammo_Hung
Sammy "The Bull" Gravano	http://en.wikipedia.org/wiki/Sammy_%22The_Bull%22_Gravano
Sammy Baugh	http://en.wikipedia.org/wiki/Sammy_Baugh
Sammy Cahn	http://en.wikipedia.org/wiki/Sammy_Cahn
Sammy Davis, Jr.	http://en.wikipedia.org/wiki/Sammy_Davis%2C_Jr.
Sammy Hagar	http://en.wikipedia.org/wiki/Sammy_Hagar
Sammy Sosa	http://en.wikipedia.org/wiki/Sammy_Sosa
Sammy Wilson	http://en.wikipedia.org/wiki/Sammy_Wilson
Samson Occom	http://en.wikipedia.org/wiki/Samson_Occom
Samuel A. Foote	http://en.wikipedia.org/wiki/Samuel_A._Foote
Samuel Adams	http://en.wikipedia.org/wiki/Samuel_Adams
Samuel Alito	http://en.wikipedia.org/wiki/Samuel_Alito
Samuel Bailey	http://en.wikipedia.org/wiki/Samuel_Bailey
Samuel Barber	http://en.wikipedia.org/wiki/Samuel_Barber
Samuel Beckett	http://en.wikipedia.org/wiki/Samuel_Beckett
Samuel Butler	http://en.wikipedia.org/wiki/Samuel_Butler_(novelist)
Samuel Butler	http://en.wikipedia.org/wiki/Samuel_Butler_(poet)
Samuel Butler	http://en.wikipedia.org/wiki/Samuel_Butler_(schoolmaster)
Samuel C. C. Ting	http://en.wikipedia.org/wiki/Samuel_C._C._Ting
Samuel Clarke	http://en.wikipedia.org/wiki/Samuel_Clarke
Samuel Colt	http://en.wikipedia.org/wiki/Samuel_Colt
Samuel Crompton	http://en.wikipedia.org/wiki/Samuel_Crompton
Samuel Crowther	http://en.wikipedia.org/wiki/Samuel_Crowther
Samuel de Champlain	http://en.wikipedia.org/wiki/Samuel_de_Champlain
Samuel Eliot Morison	http://en.wikipedia.org/wiki/Samuel_Eliot_Morison
Samuel F. B. Morse	http://en.wikipedia.org/wiki/Samuel_F._B._Morse
Samuel Foote	http://en.wikipedia.org/wiki/Samuel_Foote
Samuel Fuller	http://en.wikipedia.org/wiki/Samuel_Fuller
Samuel Goldwyn	http://en.wikipedia.org/wiki/Samuel_Goldwyn
Samuel Gompers	http://en.wikipedia.org/wiki/Samuel_Gompers
Samuel Goudsmit	http://en.wikipedia.org/wiki/Samuel_Goudsmit
Samuel Gridley Howe	http://en.wikipedia.org/wiki/Samuel_Gridley_Howe
Samuel Hahnemann	http://en.wikipedia.org/wiki/Samuel_Hahnemann
Samuel Hearne	http://en.wikipedia.org/wiki/Samuel_Hearne
Samuel Hood	http://en.wikipedia.org/wiki/Samuel_Hood,_1st_Viscount_Hood
Samuel Hopkins	http://en.wikipedia.org/wiki/Samuel_Hopkins_(1721-1803)
Samuel Hopkins Adams	http://en.wikipedia.org/wiki/Samuel_Hopkins_Adams
Samuel J. Palmisano	http://en.wikipedia.org/wiki/Samuel_J._Palmisano
Samuel J. Tilden	http://en.wikipedia.org/wiki/Samuel_J._Tilden
Samuel Jackson Randall	http://en.wikipedia.org/wiki/Samuel_Jackson_Randall
Samuel Johnson	http://en.wikipedia.org/wiki/Samuel_Johnson
Samuel K. Skinner	http://en.wikipedia.org/wiki/Samuel_K._Skinner
Samuel L. Jackson	http://en.wikipedia.org/wiki/Samuel_L._Jackson
Samuel Liddell MacGregor Mathers	http://en.wikipedia.org/wiki/Samuel_Liddell_MacGregor_Mathers
Samuel Lover	http://en.wikipedia.org/wiki/Samuel_Lover
Samuel P. Bush	http://en.wikipedia.org/wiki/Samuel_P._Bush
Samuel P. Huntington	http://en.wikipedia.org/wiki/Samuel_P._Huntington
Samuel Palmer	http://en.wikipedia.org/wiki/Samuel_Palmer
Samuel Pepys	http://en.wikipedia.org/wiki/Samuel_Pepys
Samuel R. Delany	http://en.wikipedia.org/wiki/Samuel_R._Delany
Samuel Richardson	http://en.wikipedia.org/wiki/Samuel_Richardson
Samuel S. Stratton	http://en.wikipedia.org/wiki/Samuel_S._Stratton
Samuel Taylor Coleridge	http://en.wikipedia.org/wiki/Samuel_Taylor_Coleridge
Samuel W. Yorty	http://en.wikipedia.org/wiki/Samuel_W._Yorty
Sanaa Lathan	http://en.wikipedia.org/wiki/Sanaa_Lathan
Sanath Jayasuriya	http://en.wikipedia.org/wiki/Sanath_Jayasuriya
Sander M. Levin	http://en.wikipedia.org/wiki/Sander_M._Levin
Sander Vanocur	http://en.wikipedia.org/wiki/Sander_Vanocur
Sandra Bernhard	http://en.wikipedia.org/wiki/Sandra_Bernhard
Sandra Bullock	http://en.wikipedia.org/wiki/Sandra_Bullock
Sandra Day O'Connor	http://en.wikipedia.org/wiki/Sandra_Day_O%27Connor
Sandra Dee	http://en.wikipedia.org/wiki/Sandra_Dee
Sandra Lee-Vercoe	http://en.wikipedia.org/wiki/Sandra_Lee-Vercoe
Sandra Mortham	http://en.wikipedia.org/wiki/Sandra_Mortham
Sandra Oh	http://en.wikipedia.org/wiki/Sandra_Oh
Sandra Osborne	http://en.wikipedia.org/wiki/Sandra_Osborne
Sandro Botticelli	http://en.wikipedia.org/wiki/Sandro_Botticelli
Sandy Berger	http://en.wikipedia.org/wiki/Sandy_Berger
Sandy Bull	http://en.wikipedia.org/wiki/Sandy_Bull
Sandy Dennis	http://en.wikipedia.org/wiki/Sandy_Dennis
Sandy Duncan	http://en.wikipedia.org/wiki/Sandy_Duncan
Sandy Koufax	http://en.wikipedia.org/wiki/Sandy_Koufax
Sandy Levin	http://en.wikipedia.org/wiki/Sandy_Levin
Sanford D. Bishop, Jr.	http://en.wikipedia.org/wiki/Sanford_D._Bishop%2C_Jr.
Sani Abacha	http://en.wikipedia.org/wiki/Sani_Abacha
Sania Mirza	http://en.wikipedia.org/wiki/Sania_Mirza
Sanjay Dutt	http://en.wikipedia.org/wiki/Sanjay_Dutt
Sanjay Gupta	http://en.wikipedia.org/wiki/Sanjay_Gupta
Sanjay Kumar	http://en.wikipedia.org/wiki/Sanjay_Kumar
Santiago Amigorena	http://en.wikipedia.org/wiki/Santiago_Amigorena
Santiago Calatrava	http://en.wikipedia.org/wiki/Santiago_Calatrava
Santiago Durango	http://en.wikipedia.org/wiki/Santiago_Durango
Saparmurat Niyazov	http://en.wikipedia.org/wiki/Saparmurat_Niyazov
Saparmurat Niyazov	http://en.wikipedia.org/wiki/Saparmurat_Niyazov
Sara Evans	http://en.wikipedia.org/wiki/Sara_Evans
Sara Foster	http://en.wikipedia.org/wiki/Sara_Foster
Sara Gilbert	http://en.wikipedia.org/wiki/Sara_Gilbert
Sara Paretsky	http://en.wikipedia.org/wiki/Sara_Paretsky
Sara Payson Willis Parton	http://en.wikipedia.org/wiki/Sara_Payson_Willis_Parton
Sara Rue	http://en.wikipedia.org/wiki/Sara_Rue
Sara Teasdale	http://en.wikipedia.org/wiki/Sara_Teasdale
Sarah Bernhardt	http://en.wikipedia.org/wiki/Sarah_Bernhardt
Sarah Brady	http://en.wikipedia.org/wiki/Sarah_Brady
Sarah Brightman	http://en.wikipedia.org/wiki/Sarah_Brightman
Sarah Chalke	http://en.wikipedia.org/wiki/Sarah_Chalke
Sarah Cracknell	http://en.wikipedia.org/wiki/Sarah_Cracknell
Sarah Ferguson	http://en.wikipedia.org/wiki/Sarah_Ferguson
Sarah Hughes	http://en.wikipedia.org/wiki/Sarah_Hughes
Sarah Jessica Parker	http://en.wikipedia.org/wiki/Sarah_Jessica_Parker
Sarah Josepha Hale	http://en.wikipedia.org/wiki/Sarah_Josepha_Hale
Sarah Kemble Knight	http://en.wikipedia.org/wiki/Sarah_Kemble_Knight
Sarah Marbeck	http://en.wikipedia.org/wiki/Sarah_Marbeck
Sarah McClendon	http://en.wikipedia.org/wiki/Sarah_McClendon
Sarah McLachlan	http://en.wikipedia.org/wiki/Sarah_McLachlan
Sarah Michelle Gellar	http://en.wikipedia.org/wiki/Sarah_Michelle_Gellar
Sarah Miles	http://en.wikipedia.org/wiki/Sarah_Miles
Sarah Newton	http://en.wikipedia.org/wiki/Sarah_Newton
Sarah Orne Jewett	http://en.wikipedia.org/wiki/Sarah_Orne_Jewett
Sarah Palin	http://en.wikipedia.org/wiki/Sarah_Palin
Sarah Paulson	http://en.wikipedia.org/wiki/Sarah_Paulson
Sarah Polley	http://en.wikipedia.org/wiki/Sarah_Polley
Sarah Siddons	http://en.wikipedia.org/wiki/Sarah_Siddons
Sarah Silverman	http://en.wikipedia.org/wiki/Sarah_Silverman
Sarah Susanka	http://en.wikipedia.org/wiki/Sarah_Susanka
Sarah Sutton	http://en.wikipedia.org/wiki/Sarah_Sutton
Sarah Teather	http://en.wikipedia.org/wiki/Sarah_Teather
Sarah Vaughan	http://en.wikipedia.org/wiki/Sarah_Vaughan
Sarah Vowell	http://en.wikipedia.org/wiki/Sarah_Vowell
Sarah Wentworth Morton	http://en.wikipedia.org/wiki/Sarah_Wentworth_Morton
Sarah Wollaston	http://en.wikipedia.org/wiki/Sarah_Wollaston
Sarah Zettel	http://en.wikipedia.org/wiki/Sarah_Zettel
Sargent Shriver	http://en.wikipedia.org/wiki/Sargent_Shriver
Sasha Alexander	http://en.wikipedia.org/wiki/Sasha_Alexander
Sasha Mitchell	http://en.wikipedia.org/wiki/Sasha_Mitchell
Satchel Paige	http://en.wikipedia.org/wiki/Satchel_Paige
Saul Bellow	http://en.wikipedia.org/wiki/Saul_Bellow
Saxby Chambliss	http://en.wikipedia.org/wiki/Saxby_Chambliss
Sayyid Qutb	http://en.wikipedia.org/wiki/Sayyid_Qutb
Scarlett Johansson	http://en.wikipedia.org/wiki/Scarlett_Johansson
Scatman Crothers	http://en.wikipedia.org/wiki/Scatman_Crothers
Schuyler Colfax	http://en.wikipedia.org/wiki/Schuyler_Colfax
Schuyler Fisk	http://en.wikipedia.org/wiki/Schuyler_Fisk
Scipio Africanus	http://en.wikipedia.org/wiki/Scipio_Africanus
Scooter Ward	http://en.wikipedia.org/wiki/Scooter_Ward
Scott Adams	http://en.wikipedia.org/wiki/Scott_Adams
Scott Adams	http://en.wikipedia.org/wiki/Scott_Adams_(game_designer)
Scott Adams	http://en.wikipedia.org/wiki/Scott_Adams
Scott Baio	http://en.wikipedia.org/wiki/Scott_Baio
Scott Bairstow	http://en.wikipedia.org/wiki/Scott_Bairstow
Scott Bakula	http://en.wikipedia.org/wiki/Scott_Bakula
Scott Brown	http://en.wikipedia.org/wiki/Scott_Brown
Scott C. Bone	http://en.wikipedia.org/wiki/Scott_C._Bone
Scott Caan	http://en.wikipedia.org/wiki/Scott_Caan
Scott Carpenter	http://en.wikipedia.org/wiki/Scott_Carpenter
Scott English	http://en.wikipedia.org/wiki/Scott_English
Scott Foley	http://en.wikipedia.org/wiki/Scott_Foley
Scott G. McNealy	http://en.wikipedia.org/wiki/Scott_G._McNealy
Scott Garrett	http://en.wikipedia.org/wiki/Scott_Garrett
Scott Glenn	http://en.wikipedia.org/wiki/Scott_Glenn
Scott Hamilton	http://en.wikipedia.org/wiki/Scott_Hamilton_(figure_skater)
Scott Herren	http://en.wikipedia.org/wiki/Scott_Herren
Scott Horton	http://en.wikipedia.org/wiki/Scott_Horton_(lawyer)
Scott Ian	http://en.wikipedia.org/wiki/Scott_Ian
Scott Joplin	http://en.wikipedia.org/wiki/Scott_Joplin
Scott Kirkland	http://en.wikipedia.org/wiki/Scott_Kirkland
Scott Levy	http://en.wikipedia.org/wiki/Scott_Levy_(actor)
Scott Lowell	http://en.wikipedia.org/wiki/Scott_Lowell
Scott McCallum	http://en.wikipedia.org/wiki/Scott_McCallum
Scott McClellan	http://en.wikipedia.org/wiki/Scott_McClellan
Scott McCloud	http://en.wikipedia.org/wiki/Scott_McCloud
Scott McInnis	http://en.wikipedia.org/wiki/Scott_McInnis
Scott McNealy	http://en.wikipedia.org/wiki/Scott_McNealy
Scott Murphy	http://en.wikipedia.org/wiki/Scott_Murphy
Scott Patterson	http://en.wikipedia.org/wiki/Scott_Patterson_(actor)
Scott Pelley	http://en.wikipedia.org/wiki/Scott_Pelley
Scott Peterson	http://en.wikipedia.org/wiki/Scott_Peterson
Scott Ritter	http://en.wikipedia.org/wiki/Scott_Ritter
Scott Sassa	http://en.wikipedia.org/wiki/Scott_Sassa
Scott Speedman	http://en.wikipedia.org/wiki/Scott_Speedman
Scott Stapp	http://en.wikipedia.org/wiki/Scott_Stapp
Scott Thompson	http://en.wikipedia.org/wiki/Scott_Thompson
Scott Thorson	http://en.wikipedia.org/wiki/Scott_Thorson
Scott Turow	http://en.wikipedia.org/wiki/Scott_Turow
Scott Weiland	http://en.wikipedia.org/wiki/Scott_Weiland
Scott Weinger	http://en.wikipedia.org/wiki/Scott_Weinger
Scott Wolf	http://en.wikipedia.org/wiki/Scott_Wolf
Scottie Pippen	http://en.wikipedia.org/wiki/Scottie_Pippen
Scotty Moore	http://en.wikipedia.org/wiki/Scotty_Moore
Screamin' Jay Hawkins	http://en.wikipedia.org/wiki/Screamin%27_Jay_Hawkins
Seamus Heaney	http://en.wikipedia.org/wiki/Seamus_Heaney
Sean Astin	http://en.wikipedia.org/wiki/Sean_Astin
Sean Bean	http://en.wikipedia.org/wiki/Sean_Bean
Sean Biggerstaff	http://en.wikipedia.org/wiki/Sean_Biggerstaff
Sean Booth	http://en.wikipedia.org/wiki/Sean_Booth
Sean Connery	http://en.wikipedia.org/wiki/Sean_Connery
Sean Faris	http://en.wikipedia.org/wiki/Sean_Faris
Sean Flynn	http://en.wikipedia.org/wiki/Sean_Flynn
Sean Hannity	http://en.wikipedia.org/wiki/Sean_Hannity
Sean Hayes	http://en.wikipedia.org/wiki/Sean_Hayes_(actor)
Sean Kinney	http://en.wikipedia.org/wiki/Sean_Kinney
Sean Lennon	http://en.wikipedia.org/wiki/Sean_Lennon
Se�n MacBride	http://en.wikipedia.org/wiki/Se%E1n_MacBride
Sean McClory	http://en.wikipedia.org/wiki/Sean_McClory
Sean O'Casey	http://en.wikipedia.org/wiki/Sean_O%27Casey
Sean O'Faolain	http://en.wikipedia.org/wiki/Sean_O%27Faolain
Sean Patrick Flanery	http://en.wikipedia.org/wiki/Sean_Patrick_Flanery
Sean Patrick Thomas	http://en.wikipedia.org/wiki/Sean_Patrick_Thomas
Sean Paul	http://en.wikipedia.org/wiki/Sean_Paul
Sean Penn	http://en.wikipedia.org/wiki/Sean_Penn
Sean Wilentz	http://en.wikipedia.org/wiki/Sean_Wilentz
Sean Young	http://en.wikipedia.org/wiki/Sean_Young
Seann William Scott	http://en.wikipedia.org/wiki/Seann_William_Scott
Sebastian Bach	http://en.wikipedia.org/wiki/Sebastian_Bach
Sebastian Brant	http://en.wikipedia.org/wiki/Sebastian_Brant
Sebastian Cabot	http://en.wikipedia.org/wiki/Sebastian_Cabot_(actor)
Sebastian Cabot	http://en.wikipedia.org/wiki/Sebastian_Cabot_(explorer)
Sebastian Coe	http://en.wikipedia.org/wiki/Sebastian_Coe
Sebastian Franck	http://en.wikipedia.org/wiki/Sebastian_Franck
Sebastian Junger	http://en.wikipedia.org/wiki/Sebastian_Junger
Sebasti�n Lerdo de Tejada	http://en.wikipedia.org/wiki/Sebasti%E1n_Lerdo_de_Tejada
Sebastian M�nster	http://en.wikipedia.org/wiki/Sebastian_M%FCnster
Sebasti�n Pi�era	http://en.wikipedia.org/wiki/Sebasti%E1n_Pi%F1era
S�bastien de Vauban	http://en.wikipedia.org/wiki/S%E9bastien_de_Vauban
Sela Ward	http://en.wikipedia.org/wiki/Sela_Ward
Selim I	http://en.wikipedia.org/wiki/Selim_I
Selim II	http://en.wikipedia.org/wiki/Selim_II
Sellapan Ramanathan	http://en.wikipedia.org/wiki/Sellapan_Ramanathan
Selma Blair	http://en.wikipedia.org/wiki/Selma_Blair
Selma Lagerl�f	http://en.wikipedia.org/wiki/Selma_Lagerl%F6f
Sepp Blatter	http://en.wikipedia.org/wiki/Sepp_Blatter
Sepp Dietrich	http://en.wikipedia.org/wiki/Sepp_Dietrich
Septimius Severus	http://en.wikipedia.org/wiki/Septimius_Severus
Serena Williams	http://en.wikipedia.org/wiki/Serena_Williams
Serge Clair	http://en.wikipedia.org/wiki/Serge_Clair
Serge Gainsbourg	http://en.wikipedia.org/wiki/Serge_Gainsbourg
Serge Reggiani	http://en.wikipedia.org/wiki/Serge_Reggiani
Sergei Eisenstein	http://en.wikipedia.org/wiki/Sergei_Eisenstein
Sergei Parajanov	http://en.wikipedia.org/wiki/Sergei_Parajanov
Sergei Prokofiev	http://en.wikipedia.org/wiki/Sergei_Prokofiev
Sergei Rachmaninov	http://en.wikipedia.org/wiki/Sergei_Rachmaninov
Sergei Sidorsky	http://en.wikipedia.org/wiki/Sergei_Sidorsky
Sergei Stanishev	http://en.wikipedia.org/wiki/Sergei_Stanishev
Sergei Stepashin	http://en.wikipedia.org/wiki/Sergei_Stepashin
Sergey Abramov	http://en.wikipedia.org/wiki/Sergey_Abramov
Sergey Bagapsh	http://en.wikipedia.org/wiki/Sergey_Bagapsh
Sergey Brin	http://en.wikipedia.org/wiki/Sergey_Brin
Sergey Sidorsky	http://en.wikipedia.org/wiki/Sergey_Sidorsky
Sergio Amidei	http://en.wikipedia.org/wiki/Sergio_Amidei
Sergio Aragones	http://en.wikipedia.org/wiki/Sergio_Aragones
Sergio de Mello	http://en.wikipedia.org/wiki/Sergio_de_Mello
Sergio Leone	http://en.wikipedia.org/wiki/Sergio_Leone
Sergio Mendes	http://en.wikipedia.org/wiki/Sergio_Mendes
Sergio Osme�a	http://en.wikipedia.org/wiki/Sergio_Osme%F1a
Serj Tankian	http://en.wikipedia.org/wiki/Serj_Tankian
Serphin Maltese	http://en.wikipedia.org/wiki/Serphin_Maltese
Servius Sulpicius Rufus	http://en.wikipedia.org/wiki/Servius_Sulpicius_Rufus
Serzh Sargsyan	http://en.wikipedia.org/wiki/Serzh_Sargsyan
Sessue Hayakawa	http://en.wikipedia.org/wiki/Sessue_Hayakawa
Sete Gibernau	http://en.wikipedia.org/wiki/Sete_Gibernau
Seth Green	http://en.wikipedia.org/wiki/Seth_Green
Seth MacFarlane	http://en.wikipedia.org/wiki/Seth_MacFarlane
Seth Meyers	http://en.wikipedia.org/wiki/Seth_Meyers
Severiano Ballesteros	http://en.wikipedia.org/wiki/Severiano_Ballesteros
Severina Vuckovic	http://en.wikipedia.org/wiki/Severina_Vuckovic
Severo Sarduy	http://en.wikipedia.org/wiki/Severo_Sarduy
Severus Alexander	http://en.wikipedia.org/wiki/Severus_Alexander
Sewall Wright	http://en.wikipedia.org/wiki/Sewall_Wright
Seymour Cray	http://en.wikipedia.org/wiki/Seymour_Cray
Seymour Hersh	http://en.wikipedia.org/wiki/Seymour_Hersh
Seymour Papert	http://en.wikipedia.org/wiki/Seymour_Papert
Shabana Mahmood	http://en.wikipedia.org/wiki/Shabana_Mahmood
Shabba Ranks	http://en.wikipedia.org/wiki/Shabba_Ranks
Shadoe Stevens	http://en.wikipedia.org/wiki/Shadoe_Stevens
Shaggy 2 Dope	http://en.wikipedia.org/wiki/Shaggy_2_Dope
Shah of Iran	http://en.wikipedia.org/wiki/Mohammed_Reza_Pahlavi
Shahid Afridi	http://en.wikipedia.org/wiki/Shahid_Afridi
Shahrukh Khan	http://en.wikipedia.org/wiki/Shahrukh_Khan
Shailesh Vara	http://en.wikipedia.org/wiki/Shailesh_Vara
Shaka Zulu	http://en.wikipedia.org/wiki/Shaka_Zulu
Shakin' Stevens	http://en.wikipedia.org/wiki/Shakin%27_Stevens
Shalom Harlow	http://en.wikipedia.org/wiki/Shalom_Harlow
Shamsi Vuai Nahodha	http://en.wikipedia.org/wiki/Shamsi_Vuai_Nahodha
Shana Alexander	http://en.wikipedia.org/wiki/Shana_Alexander
Shane Barbi	http://en.wikipedia.org/wiki/Shane_Barbi
Shane MacGowan	http://en.wikipedia.org/wiki/Shane_MacGowan
Shane Warne	http://en.wikipedia.org/wiki/Shane_Warne
Shane West	http://en.wikipedia.org/wiki/Shane_West
Shania Twain	http://en.wikipedia.org/wiki/Shania_Twain
Shannen Doherty	http://en.wikipedia.org/wiki/Shannen_Doherty
Shannon Elizabeth	http://en.wikipedia.org/wiki/Shannon_Elizabeth
Shannon Hoon	http://en.wikipedia.org/wiki/Shannon_Hoon
Shannon Lee	http://en.wikipedia.org/wiki/Shannon_Lee
Shannon Lucid	http://en.wikipedia.org/wiki/Shannon_Lucid
Shannyn Sossamon	http://en.wikipedia.org/wiki/Shannyn_Sossamon
Shapur I	http://en.wikipedia.org/wiki/Shapur_I
Shapur II	http://en.wikipedia.org/wiki/Shapur_II
Shaquille O'Neal	http://en.wikipedia.org/wiki/Shaquille_O%27Neal
Shar Jackson	http://en.wikipedia.org/wiki/Shar_Jackson
Shari Belafonte	http://en.wikipedia.org/wiki/Shari_Belafonte
Shari Lewis	http://en.wikipedia.org/wiki/Shari_Lewis
Sharif Ahmed	http://en.wikipedia.org/wiki/Sharif_Ahmed
Sharon Gless	http://en.wikipedia.org/wiki/Sharon_Gless
Sharon Hodgson	http://en.wikipedia.org/wiki/Sharon_Hodgson
Sharon Lawrence	http://en.wikipedia.org/wiki/Sharon_Lawrence
Sharon Leal	http://en.wikipedia.org/wiki/Sharon_Leal
Sharon Olds	http://en.wikipedia.org/wiki/Sharon_Olds
Sharon Osbourne	http://en.wikipedia.org/wiki/Sharon_Osbourne
Sharon Stone	http://en.wikipedia.org/wiki/Sharon_Stone
Sharon Tate	http://en.wikipedia.org/wiki/Sharon_Tate
Shaukat Aziz	http://en.wikipedia.org/wiki/Shaukat_Aziz
Shaukat Aziz	http://en.wikipedia.org/wiki/Shaukat_Aziz
Shaun Cassidy	http://en.wikipedia.org/wiki/Shaun_Cassidy
Shaun Donovan	http://en.wikipedia.org/wiki/Shaun_Donovan
Shaun Pollock	http://en.wikipedia.org/wiki/Shaun_Pollock
Shaun White	http://en.wikipedia.org/wiki/Shaun_White
Shaun Woodward	http://en.wikipedia.org/wiki/Shaun_Woodward
Shavkat Mirziyayev	http://en.wikipedia.org/wiki/Shavkat_Mirziyayev
Shawn Ashmore	http://en.wikipedia.org/wiki/Shawn_Ashmore
Shawn Colvin	http://en.wikipedia.org/wiki/Shawn_Colvin
Shawn Fanning	http://en.wikipedia.org/wiki/Shawn_Fanning
Shawn Levy	http://en.wikipedia.org/wiki/Shawn_Anthony_Levy
Shawn Michaels	http://en.wikipedia.org/wiki/Shawn_Michaels
Shawn Wayans	http://en.wikipedia.org/wiki/Shawn_Wayans
Shawnee Smith	http://en.wikipedia.org/wiki/Shawnee_Smith
Sheb Wooley	http://en.wikipedia.org/wiki/Sheb_Wooley
Shecky Greene	http://en.wikipedia.org/wiki/Shecky_Greene
Sheena Easton	http://en.wikipedia.org/wiki/Sheena_Easton
Sheeri Rappaport	http://en.wikipedia.org/wiki/Sheeri_Rappaport
Sheik Hamad bin Khalifa al-Thani	http://en.wikipedia.org/wiki/Hamad_bin_Khalifa_Al_Thani
Sheikh Ahmed Yassin	http://en.wikipedia.org/wiki/Sheikh_Ahmed_Yassin
Sheikh Hasina	http://en.wikipedia.org/wiki/Sheikh_Hasina
Sheila E	http://en.wikipedia.org/wiki/Sheila_E
Sheila Gilmore	http://en.wikipedia.org/wiki/Sheila_Gilmore
Sheila Hancock	http://en.wikipedia.org/wiki/Sheila_Hancock
Sheila Jackson Lee	http://en.wikipedia.org/wiki/Sheila_Jackson_Lee
Sheila Kaye-Smith	http://en.wikipedia.org/wiki/Sheila_Kaye-Smith
Sheila Kuehl	http://en.wikipedia.org/wiki/Sheila_Kuehl
Sheilah Graham	http://en.wikipedia.org/wiki/Sheilah_Graham
Shel Silverstein	http://en.wikipedia.org/wiki/Shel_Silverstein
Shelby Foote	http://en.wikipedia.org/wiki/Shelby_Foote
Shelby Lynne	http://en.wikipedia.org/wiki/Shelby_Lynne
Shelby Steele	http://en.wikipedia.org/wiki/Shelby_Steele
Sheldon Adelson	http://en.wikipedia.org/wiki/Sheldon_Adelson
Sheldon Glashow	http://en.wikipedia.org/wiki/Sheldon_Glashow
Sheldon Whitehouse	http://en.wikipedia.org/wiki/Sheldon_Whitehouse
Shelley Berkley	http://en.wikipedia.org/wiki/Shelley_Berkley
Shelley Duvall	http://en.wikipedia.org/wiki/Shelley_Duvall
Shelley Fabares	http://en.wikipedia.org/wiki/Shelley_Fabares
Shelley Hack	http://en.wikipedia.org/wiki/Shelley_Hack
Shelley Long	http://en.wikipedia.org/wiki/Shelley_Long
Shelley Malil	http://en.wikipedia.org/wiki/Shelley_Malil
Shelley Moore Capito	http://en.wikipedia.org/wiki/Shelley_Moore_Capito
Shelley Morrison	http://en.wikipedia.org/wiki/Shelley_Morrison
Shelley Winters	http://en.wikipedia.org/wiki/Shelley_Winters
Shemar Moore	http://en.wikipedia.org/wiki/Shemar_Moore
Shemp Howard	http://en.wikipedia.org/wiki/Shemp_Howard
Shepard Smith	http://en.wikipedia.org/wiki/Shepard_Smith
Shere Hite	http://en.wikipedia.org/wiki/Shere_Hite
Sheree North	http://en.wikipedia.org/wiki/Sheree_North
Sheri S. Tepper	http://en.wikipedia.org/wiki/Sheri_S._Tepper
Sherilyn Fenn	http://en.wikipedia.org/wiki/Sherilyn_Fenn
Sherman Adams	http://en.wikipedia.org/wiki/Sherman_Adams
Sherman Alexie	http://en.wikipedia.org/wiki/Sherman_Alexie
Sherman Austin	http://en.wikipedia.org/wiki/Sherman_Austin
Sherman Hemsley	http://en.wikipedia.org/wiki/Sherman_Hemsley
Sherman W. Tribbitt	http://en.wikipedia.org/wiki/Sherman_W._Tribbitt
Sherrod Brown	http://en.wikipedia.org/wiki/Sherrod_Brown
Sherry Alberoni	http://en.wikipedia.org/wiki/Sherry_Alberoni
Sherry Lansing	http://en.wikipedia.org/wiki/Sherry_Lansing
Sherry Stringfield	http://en.wikipedia.org/wiki/Sherry_Stringfield
Sherwood Anderson	http://en.wikipedia.org/wiki/Sherwood_Anderson
Sherwood Boehlert	http://en.wikipedia.org/wiki/Sherwood_Boehlert
Sherwood Boehlert	http://en.wikipedia.org/wiki/Sherwood_Boehlert
Sherwood Schwartz	http://en.wikipedia.org/wiki/Sherwood_Schwartz
Sheryl Crow	http://en.wikipedia.org/wiki/Sheryl_Crow
Sheryl Lee	http://en.wikipedia.org/wiki/Sheryl_Lee
Sheryl Swoopes	http://en.wikipedia.org/wiki/Sheryl_Swoopes
Sheryll Murray	http://en.wikipedia.org/wiki/Sheryll_Murray
Shia LaBeouf	http://en.wikipedia.org/wiki/Shia_LaBeouf
Shigeru Miyamoto	http://en.wikipedia.org/wiki/Shigeru_Miyamoto
Shigeru Yoshida	http://en.wikipedia.org/wiki/Shigeru_Yoshida
Shimon Peres	http://en.wikipedia.org/wiki/Shimon_Peres
Shin Amano	http://en.wikipedia.org/wiki/Shin_Amano
Shiri Appleby	http://en.wikipedia.org/wiki/Shiri_Appleby
Shirin Ebadi	http://en.wikipedia.org/wiki/Shirin_Ebadi
Shirley A. Jackson	http://en.wikipedia.org/wiki/Shirley_Jackson_(physicist)
Shirley Ann Grau	http://en.wikipedia.org/wiki/Shirley_Ann_Grau
Shirley Bassey	http://en.wikipedia.org/wiki/Shirley_Bassey
Shirley Booth	http://en.wikipedia.org/wiki/Shirley_Booth
Shirley Chisholm	http://en.wikipedia.org/wiki/Shirley_Chisholm
Shirley Franklin	http://en.wikipedia.org/wiki/Shirley_Franklin
Shirley Hazzard	http://en.wikipedia.org/wiki/Shirley_Hazzard
Shirley Horn	http://en.wikipedia.org/wiki/Shirley_Horn
Shirley Hughes	http://en.wikipedia.org/wiki/Shirley_Hughes
Shirley Jackson	http://en.wikipedia.org/wiki/Shirley_Jackson
Shirley Jones	http://en.wikipedia.org/wiki/Shirley_Jones
Shirley M. Tilghman	http://en.wikipedia.org/wiki/Shirley_M._Tilghman
Shirley MacLaine	http://en.wikipedia.org/wiki/Shirley_MacLaine
Shirley Manson	http://en.wikipedia.org/wiki/Shirley_Manson
Shirley Temple	http://en.wikipedia.org/wiki/Shirley_Temple
Shoaib Akhtar	http://en.wikipedia.org/wiki/Shoaib_Akhtar
Shock G	http://en.wikipedia.org/wiki/Shock_G
Shoeless Joe Jackson	http://en.wikipedia.org/wiki/Shoeless_Joe_Jackson
Shoko Asahara	http://en.wikipedia.org/wiki/Shoko_Asahara
Sholem Asch	http://en.wikipedia.org/wiki/Sholem_Asch
Shooby Taylor	http://en.wikipedia.org/wiki/Shooby_Taylor
Shukri Ghanem	http://en.wikipedia.org/wiki/Shukri_Ghanem
Sia Barbi	http://en.wikipedia.org/wiki/Sia_Barbi
Si�n C. James	http://en.wikipedia.org/wiki/Sian_James_(politician)
Sibel Edmonds	http://en.wikipedia.org/wiki/Sibel_Edmonds
Sid Caesar	http://en.wikipedia.org/wiki/Sid_Caesar
Sid James	http://en.wikipedia.org/wiki/Sid_James
Sid Krofft	http://en.wikipedia.org/wiki/Sid_Krofft
Sid Meier	http://en.wikipedia.org/wiki/Sid_Meier
Sid Morrison	http://en.wikipedia.org/wiki/Sid_Morrison
Sid Vicious	http://en.wikipedia.org/wiki/Sid_Vicious
Sidi Mohamed Ould Boubacar	http://en.wikipedia.org/wiki/Sidi_Mohamed_Ould_Boubacar
Sidney Altman	http://en.wikipedia.org/wiki/Sidney_Altman
Sidney Blackmer	http://en.wikipedia.org/wiki/Sidney_Blackmer
Sidney Blumenthal	http://en.wikipedia.org/wiki/Sidney_Blumenthal
Sidney Coe Howard	http://en.wikipedia.org/wiki/Sidney_Coe_Howard
Sidney D. Drell	http://en.wikipedia.org/wiki/Sidney_D._Drell
Sidney Hook	http://en.wikipedia.org/wiki/Sidney_Hook
Sidney J. Furie	http://en.wikipedia.org/wiki/Sidney_J._Furie
Sidney Lanfield	http://en.wikipedia.org/wiki/Sidney_Lanfield
Sidney Lanier	http://en.wikipedia.org/wiki/Sidney_Lanier
Sidney Lumet	http://en.wikipedia.org/wiki/Sidney_Lumet
Sidney Poitier	http://en.wikipedia.org/wiki/Sidney_Poitier
Sidney R. Yates	http://en.wikipedia.org/wiki/Sidney_R._Yates
Sidney Sheldon	http://en.wikipedia.org/wiki/Sidney_Sheldon
Sidney Souers	http://en.wikipedia.org/wiki/Sidney_Souers
Siegfried Fischbacher	http://en.wikipedia.org/wiki/Siegfried_Fischbacher
Siegfried Sassoon	http://en.wikipedia.org/wiki/Siegfried_Sassoon
Sienna Guillory	http://en.wikipedia.org/wiki/Sienna_Guillory
Sienna Miller	http://en.wikipedia.org/wiki/Sienna_Miller
Sigismond Thalberg	http://en.wikipedia.org/wiki/Sigismond_Thalberg
Sigmund Freud	http://en.wikipedia.org/wiki/Sigmund_Freud
Signe Hasso	http://en.wikipedia.org/wiki/Signe_Hasso
Sigourney Weaver	http://en.wikipedia.org/wiki/Sigourney_Weaver
Sigtryggur Baldursson	http://en.wikipedia.org/wiki/Sigtryggur_Baldursson
Siim Kallas	http://en.wikipedia.org/wiki/Siim_Kallas
Sila Calder�n	http://en.wikipedia.org/wiki/Sila_Calder%F3n
Silas Deane	http://en.wikipedia.org/wiki/Silas_Deane
Silas Wright	http://en.wikipedia.org/wiki/Silas_Wright
Silkk the Shocker	http://en.wikipedia.org/wiki/Silkk_the_Shocker
Silvan Shalom	http://en.wikipedia.org/wiki/Silvan_Shalom
Silvana Mangano	http://en.wikipedia.org/wiki/Silvana_Mangano
Silvestre Reyes	http://en.wikipedia.org/wiki/Silvestre_Reyes
Silvio Amadio	http://en.wikipedia.org/wiki/Silvio_Amadio
Silvio Berlusconi	http://en.wikipedia.org/wiki/Silvio_Berlusconi
Silvio O. Conte	http://en.wikipedia.org/wiki/Silvio_O._Conte
Silvio Pellico	http://en.wikipedia.org/wiki/Silvio_Pellico
Sim�on-Denis Poisson	http://en.wikipedia.org/wiki/Sim%E9on-Denis_Poisson
Simon Abkarian	http://en.wikipedia.org/wiki/Simon_Abkarian
Simon Baker	http://en.wikipedia.org/wiki/Simon_Baker
Simon ben Yohai	http://en.wikipedia.org/wiki/Simon_ben_Yohai
Sim�n Bol�var	http://en.wikipedia.org/wiki/Sim%F3n_Bol%EDvar
Simon Burns	http://en.wikipedia.org/wiki/Simon_Burns
Simon Callow	http://en.wikipedia.org/wiki/Simon_Callow
Simon Conway Morris	http://en.wikipedia.org/wiki/Simon_Conway_Morris
Simon Cowell	http://en.wikipedia.org/wiki/Simon_Cowell
Simon Dach	http://en.wikipedia.org/wiki/Simon_Dach
Simon Danczuk	http://en.wikipedia.org/wiki/Simon_Danczuk
Simon Hart	http://en.wikipedia.org/wiki/Simon_Hart
Simon Hughes	http://en.wikipedia.org/wiki/Simon_Hughes
Simon Kirby	http://en.wikipedia.org/wiki/Simon_Kirby
Simon Kuznets	http://en.wikipedia.org/wiki/Simon_Kuznets
Simon Le Bon	http://en.wikipedia.org/wiki/Simon_Le_Bon
Simon Mills	http://en.wikipedia.org/wiki/Simon_Mills
Simon Newcomb	http://en.wikipedia.org/wiki/Simon_Newcomb
Simon of Sudbury	http://en.wikipedia.org/wiki/Simon_of_Sudbury
Simon Pegg	http://en.wikipedia.org/wiki/Simon_Pegg
Simon Raymonde	http://en.wikipedia.org/wiki/Simon_Raymonde
Simon Reevell	http://en.wikipedia.org/wiki/Simon_Reevell
Simon Rex	http://en.wikipedia.org/wiki/Simon_Rex
Simon Stevin	http://en.wikipedia.org/wiki/Simon_Stevin
Simon van der Meer	http://en.wikipedia.org/wiki/Simon_van_der_Meer
Simon Wiesenthal	http://en.wikipedia.org/wiki/Simon_Wiesenthal
Simon Winchester	http://en.wikipedia.org/wiki/Simon_Winchester
Simon Wright	http://en.wikipedia.org/wiki/Simon_Wright_(politician)
Simone de Beauvoir	http://en.wikipedia.org/wiki/Simone_de_Beauvoir
Simone Martini	http://en.wikipedia.org/wiki/Simone_Martini
Simone Signoret	http://en.wikipedia.org/wiki/Simone_Signoret
Simone Simon	http://en.wikipedia.org/wiki/Simone_Simon
Simonides of Amorgos	http://en.wikipedia.org/wiki/Simonides_of_Amorgos
Simonides of Ceos	http://en.wikipedia.org/wiki/Simonides_of_Ceos
Sinclair Lewis	http://en.wikipedia.org/wiki/Sinclair_Lewis
Sinclair Ross	http://en.wikipedia.org/wiki/Sinclair_Ross
Sin�ad Cusack	http://en.wikipedia.org/wiki/Sin%E9ad_Cusack
Sinead O'Connor	http://en.wikipedia.org/wiki/Sinead_O%27Connor
Sin-Itiro Tomonaga	http://en.wikipedia.org/wiki/Sin-Itiro_Tomonaga
Siobhain McDonagh	http://en.wikipedia.org/wiki/Siobhain_McDonagh
Siobhan Fahey	http://en.wikipedia.org/wiki/Siobhan_Fahey
Siouxsie Sioux	http://en.wikipedia.org/wiki/Siouxsie_Sioux
Sir Alex Ferguson	http://en.wikipedia.org/wiki/Sir_Alex_Ferguson
Sir Alf Ramsey	http://en.wikipedia.org/wiki/Sir_Alf_Ramsey
Sir Allan Kemakeza	http://en.wikipedia.org/wiki/Sir_Allan_Kemakeza
Sir Anerood Jugnauth	http://en.wikipedia.org/wiki/Sir_Anerood_Jugnauth
Sir Anthony Panizzi	http://en.wikipedia.org/wiki/Sir_Anthony_Panizzi
Sir Anthony Shirley	http://en.wikipedia.org/wiki/Sir_Anthony_Shirley
Sir Banastre Tarleton	http://en.wikipedia.org/wiki/Sir_Banastre_Tarleton
Sir Benjamin Baker	http://en.wikipedia.org/wiki/Sir_Benjamin_Baker
Sir Bobby Robson	http://en.wikipedia.org/wiki/Sir_Bobby_Robson
Sir Charles Bell	http://en.wikipedia.org/wiki/Sir_Charles_Bell
Sir Charles G. D. Roberts	http://en.wikipedia.org/wiki/Sir_Charles_G._D._Roberts
Sir Charles Hall�	http://en.wikipedia.org/wiki/Sir_Charles_Hall%E9
Sir Christopher Hatton	http://en.wikipedia.org/wiki/Sir_Christopher_Hatton
Sir Clifford Husbands	http://en.wikipedia.org/wiki/Clifford_Husbands
Sir Colville Young	http://en.wikipedia.org/wiki/Colville_Young
Sir Cuthbert Sebastian	http://en.wikipedia.org/wiki/Cuthbert_Sebastian
Sir Cyril Hinshelwood	http://en.wikipedia.org/wiki/Sir_Cyril_Hinshelwood
Sir Daniel Williams	http://en.wikipedia.org/wiki/Daniel_Williams_(Governor-General)
Sir Edward Hughes	http://en.wikipedia.org/wiki/Sir_Edward_Hughes
Sir Edward Poynter	http://en.wikipedia.org/wiki/Sir_Edward_Poynter
Sir Eyre Coote	http://en.wikipedia.org/wiki/Eyre_Coote_(East_India_Company_officer)
Sir Fabian Malbon	http://en.wikipedia.org/wiki/Sir_Fabian_Malbon
Sir Francis Drake	http://en.wikipedia.org/wiki/Sir_Francis_Drake
Sir Francis Richards	http://en.wikipedia.org/wiki/Sir_Francis_Richards
Sir Francis Walsingham	http://en.wikipedia.org/wiki/Sir_Francis_Walsingham
Sir Frederick Ballantyne	http://en.wikipedia.org/wiki/Frederick_Ballantyne
Sir Hans Sloane	http://en.wikipedia.org/wiki/Sir_Hans_Sloane
Sir Harold Kroto	http://en.wikipedia.org/wiki/Sir_Harold_Kroto
Sir Henry Bulwer	http://en.wikipedia.org/wiki/Henry_Ernest_Gascoyne_Bulwer
Sir Henry Clinton	http://en.wikipedia.org/wiki/Henry_Clinton_(American_War_of_Independence)
Sir Henry Havelock	http://en.wikipedia.org/wiki/Sir_Henry_Havelock
Sir Henry Irving	http://en.wikipedia.org/wiki/Sir_Henry_Irving
Sir Henry Parkes	http://en.wikipedia.org/wiki/Sir_Henry_Parkes
Sir Henry Percy	http://en.wikipedia.org/wiki/Henry_'Hotspur'_Percy
Sir Henry Sidney	http://en.wikipedia.org/wiki/Sir_Henry_Sidney
Sir Henry Tate	http://en.wikipedia.org/wiki/Sir_Henry_Tate
Sir Hiram Maxim	http://en.wikipedia.org/wiki/Sir_Hiram_Maxim
Sir Howard Cooke	http://en.wikipedia.org/wiki/Howard_Cooke
Sir Hudson Lowe	http://en.wikipedia.org/wiki/Hudson_Lowe
Sir Isaac Newton	http://en.wikipedia.org/wiki/Sir_Isaac_Newton
Sir Isaac Pitman	http://en.wikipedia.org/wiki/Sir_Isaac_Pitman
Sir James Carlisle	http://en.wikipedia.org/wiki/Sir_James_Carlisle
Sir James Frazer	http://en.wikipedia.org/wiki/Sir_James_Frazer
Sir James Ivory	http://en.wikipedia.org/wiki/James_Ivory_(mathematician)
Sir James Outram	http://en.wikipedia.org/wiki/Sir_James_Outram
Sir James Paget	http://en.wikipedia.org/wiki/Sir_James_Paget
Sir John Bowring	http://en.wikipedia.org/wiki/Sir_John_Bowring
Sir John Cheshire	http://en.wikipedia.org/wiki/John_Cheshire
Sir John Davies	http://en.wikipedia.org/wiki/Sir_John_Davies
Sir John Denham	http://en.wikipedia.org/wiki/Sir_John_Denham
Sir John Harington	http://en.wikipedia.org/wiki/John_Harington_(writer)
Sir John Hawkins	http://en.wikipedia.org/wiki/John_Hawkins_(author)
Sir John Hotham	http://en.wikipedia.org/wiki/Sir_John_Hotham
Sir John Oldcastle	http://en.wikipedia.org/wiki/John_Oldcastle
Sir John Scarlett	http://en.wikipedia.org/wiki/John_Scarlett
Sir John Suckling	http://en.wikipedia.org/wiki/John_Suckling_(poet)
Sir John Tenniel	http://en.wikipedia.org/wiki/Sir_John_Tenniel
Sir Joseph Banks	http://en.wikipedia.org/wiki/Sir_Joseph_Banks
Sir Leslie Stephen	http://en.wikipedia.org/wiki/Sir_Leslie_Stephen
Sir Matt Busby	http://en.wikipedia.org/wiki/Sir_Matt_Busby
Sir Matthew Hale	http://en.wikipedia.org/wiki/Sir_Matthew_Hale
Sir Michael Somare	http://en.wikipedia.org/wiki/Sir_Michael_Somare
Sir Mix-A-Lot	http://en.wikipedia.org/wiki/Sir_Mix-A-Lot
Sir Paul Haddacks	http://en.wikipedia.org/wiki/Sir_Paul_Haddacks
Sir Paulias Matane	http://en.wikipedia.org/wiki/Sir_Paulias_Matane
Sir Philip Sidney	http://en.wikipedia.org/wiki/Sir_Philip_Sidney
Sir Raymond Firth	http://en.wikipedia.org/wiki/Sir_Raymond_Firth
Sir Redvers Henry Buller	http://en.wikipedia.org/wiki/Redvers_Buller
Sir Richard Baker	http://en.wikipedia.org/wiki/Richard_Baker_(chronicler)
Sir Richard Burton	http://en.wikipedia.org/wiki/Sir_Richard_Burton
Sir Richard Empson	http://en.wikipedia.org/wiki/Sir_Richard_Empson
Sir Richard Grenville	http://en.wikipedia.org/wiki/Sir_Richard_Grenville
Sir Richard Hawkins	http://en.wikipedia.org/wiki/Sir_Richard_Hawkins
Sir Richard Owen	http://en.wikipedia.org/wiki/Sir_Richard_Owen
Sir Richard Wallace	http://en.wikipedia.org/wiki/Sir_Richard_Wallace
Sir Robert Howard	http://en.wikipedia.org/wiki/Robert_Howard_(playwright)
Sir Robert Rich	http://en.wikipedia.org/wiki/Robert_Rich,_2nd_Earl_of_Warwick
Sir Robert Robinson	http://en.wikipedia.org/wiki/Sir_Robert_Robinson
Sir Robert Sibbald	http://en.wikipedia.org/wiki/Robert_Sibbald
Sir Roger Newdigate	http://en.wikipedia.org/wiki/Sir_Roger_Newdigate
Sir Samuel Cunard	http://en.wikipedia.org/wiki/Sir_Samuel_Cunard
Sir Samuel White Baker	http://en.wikipedia.org/wiki/Sir_Samuel_White_Baker
Sir Simonds D'Ewes	http://en.wikipedia.org/wiki/Sir_Simonds_D%27Ewes
Sir Spencer Walpole	http://en.wikipedia.org/wiki/Sir_Spencer_Walpole
Sir Stamford Raffles	http://en.wikipedia.org/wiki/Sir_Stamford_Raffles
Sir Thomas Browne	http://en.wikipedia.org/wiki/Sir_Thomas_Browne
Sir Thomas Elyot	http://en.wikipedia.org/wiki/Sir_Thomas_Elyot
Sir Thomas Francis Wade	http://en.wikipedia.org/wiki/Thomas_Francis_Wade
Sir Thomas Gresham	http://en.wikipedia.org/wiki/Sir_Thomas_Gresham
Sir Thomas Lawrence	http://en.wikipedia.org/wiki/Sir_Thomas_Lawrence
Sir Thomas Lucy	http://en.wikipedia.org/wiki/Thomas_Lucy
Sir Thomas Malory	http://en.wikipedia.org/wiki/Sir_Thomas_Malory
Sir Thomas More	http://en.wikipedia.org/wiki/Sir_Thomas_More
Sir Thomas Overbury	http://en.wikipedia.org/wiki/Sir_Thomas_Overbury
Sir Thomas Wyat	http://en.wikipedia.org/wiki/Sir_Thomas_Wyat
Sir Walter Besant	http://en.wikipedia.org/wiki/Sir_Walter_Besant
Sir Walter Raleigh	http://en.wikipedia.org/wiki/Sir_Walter_Raleigh
Sir Walter Scott	http://en.wikipedia.org/wiki/Sir_Walter_Scott
Sir William Chambers	http://en.wikipedia.org/wiki/Sir_William_Chambers
Sir William Crookes	http://en.wikipedia.org/wiki/Sir_William_Crookes
Sir William Cubitt	http://en.wikipedia.org/wiki/Sir_William_Cubitt
Sir William Davenant	http://en.wikipedia.org/wiki/Sir_William_Davenant
Sir William Ramsay	http://en.wikipedia.org/wiki/Sir_William_Ramsay
Sir William Rowan Hamilton	http://en.wikipedia.org/wiki/Sir_William_Rowan_Hamilton
Sir William Temple	http://en.wikipedia.org/wiki/Sir_William_Temple
Sirhan Sirhan	http://en.wikipedia.org/wiki/Sirhan_Sirhan
Sirimavo Bandaranaike	http://en.wikipedia.org/wiki/Sirimavo_Bandaranaike
Sissy Spacek	http://en.wikipedia.org/wiki/Sissy_Spacek
Sitting Bull	http://en.wikipedia.org/wiki/Sitting_Bull
Skeet Ulrich	http://en.wikipedia.org/wiki/Skeet_Ulrich
Skeeter Davis	http://en.wikipedia.org/wiki/Skeeter_Davis
Skip Homeier	http://en.wikipedia.org/wiki/Skip_Homeier
Skip James	http://en.wikipedia.org/wiki/Skip_James
Skip Spence	http://en.wikipedia.org/wiki/Skip_Spence
Skitch Henderson	http://en.wikipedia.org/wiki/Skitch_Henderson
Slade Gorton	http://en.wikipedia.org/wiki/Slade_Gorton
Slade Gorton	http://en.wikipedia.org/wiki/Slade_Gorton
Slappy White	http://en.wikipedia.org/wiki/Slappy_White
Slick Rick	http://en.wikipedia.org/wiki/Slick_Rick
Slim Gaillard	http://en.wikipedia.org/wiki/Slim_Gaillard
Slim Jim Phantom	http://en.wikipedia.org/wiki/Slim_Jim_Phantom
Slim Pickens	http://en.wikipedia.org/wiki/Slim_Pickens
Slim Summerville	http://en.wikipedia.org/wiki/Slim_Summerville
Slim Thug	http://en.wikipedia.org/wiki/Slim_Thug
Slim Whitman	http://en.wikipedia.org/wiki/Slim_Whitman
Slobodan Milosevic	http://en.wikipedia.org/wiki/Slobodan_Milosevic
Sly Stone	http://en.wikipedia.org/wiki/Sly_Stone
Smarty Jones	http://en.wikipedia.org/wiki/Smarty_Jones
Smedley Butler	http://en.wikipedia.org/wiki/Smedley_Butler
Smokey Hormel	http://en.wikipedia.org/wiki/Smokey_Hormel
Smokey Robinson	http://en.wikipedia.org/wiki/Smokey_Robinson
Snoop Dogg	http://en.wikipedia.org/wiki/Snoop_Dogg
Snyder Rini	http://en.wikipedia.org/wiki/Snyder_Rini
Sofia Coppola	http://en.wikipedia.org/wiki/Sofia_Coppola
Sofia Vergara	http://en.wikipedia.org/wiki/Sofia_Vergara
Sojourner Truth	http://en.wikipedia.org/wiki/Sojourner_Truth
Sol Linowitz	http://en.wikipedia.org/wiki/Sol_Linowitz
Solange Knowles	http://en.wikipedia.org/wiki/Solange_Knowles
Soledad Miranda	http://en.wikipedia.org/wiki/Soledad_Miranda
Soledad O'Brien	http://en.wikipedia.org/wiki/Soledad_O%27Brien
Soleil Moon Frye	http://en.wikipedia.org/wiki/Soleil_Moon_Frye
Solomon Burke	http://en.wikipedia.org/wiki/Solomon_Burke
Solomon Linda	http://en.wikipedia.org/wiki/Solomon_Linda
Solomon Ortiz	http://en.wikipedia.org/wiki/Solomon_Ortiz
Solomon P. Ortiz	http://en.wikipedia.org/wiki/Solomon_P._Ortiz
Solomon Passy	http://en.wikipedia.org/wiki/Solomon_Passy
Solomon Zeitlin	http://en.wikipedia.org/wiki/Solomon_Zeitlin
Sonali Kulkarni	http://en.wikipedia.org/wiki/Sonali_Kulkarni
Sondra Locke	http://en.wikipedia.org/wiki/Sondra_Locke
Sonia Braga	http://en.wikipedia.org/wiki/Sonia_Braga
Sonia Gandhi	http://en.wikipedia.org/wiki/Sonia_Gandhi
Sonja Henie	http://en.wikipedia.org/wiki/Sonja_Henie
Sonny Barger	http://en.wikipedia.org/wiki/Sonny_Barger
Sonny Bono	http://en.wikipedia.org/wiki/Sonny_Bono
Sonny Callahan	http://en.wikipedia.org/wiki/Sonny_Callahan
Sonny Chiba	http://en.wikipedia.org/wiki/Sonny_Chiba
Sonny Landham	http://en.wikipedia.org/wiki/Sonny_Landham
Sonny Liston	http://en.wikipedia.org/wiki/Sonny_Liston
Sonny Montgomery	http://en.wikipedia.org/wiki/Sonny_Montgomery
Sonny Perdue	http://en.wikipedia.org/wiki/Sonny_Perdue
Sonny Perdue	http://en.wikipedia.org/wiki/Sonny_Perdue
Sonny Rollins	http://en.wikipedia.org/wiki/Sonny_Rollins
Sonny Shroyer	http://en.wikipedia.org/wiki/Sonny_Shroyer
Sonny Tufts	http://en.wikipedia.org/wiki/Sonny_Tufts
Soon-Tek Oh	http://en.wikipedia.org/wiki/Soon-Tek_Oh
Soon-Yi Previn	http://en.wikipedia.org/wiki/Soon-Yi_Previn
Sophia Bush	http://en.wikipedia.org/wiki/Sophia_Bush
Sophia Loren	http://en.wikipedia.org/wiki/Sophia_Loren
Sophie Kerr	http://en.wikipedia.org/wiki/Sophie_Kerr
Sophie Kinsella	http://en.wikipedia.org/wiki/Sophie_Kinsella
Sophie Marceau	http://en.wikipedia.org/wiki/Sophie_Marceau
S�ren Jessen-Petersen	http://en.wikipedia.org/wiki/S%F8ren_Jessen-Petersen
S�ren Kierkegaard	http://en.wikipedia.org/wiki/S%F8ren_Kierkegaard
Sorley Maclean	http://en.wikipedia.org/wiki/Sorley_Maclean
Sorrell Booke	http://en.wikipedia.org/wiki/Sorrell_Booke
Souleymane Nd�n� Ndiaye	http://en.wikipedia.org/wiki/Souleymane_Nd%E9n%E9_Ndiaye
Soupy Sales	http://en.wikipedia.org/wiki/Soupy_Sales
Sourav Ganguly	http://en.wikipedia.org/wiki/Sourav_Ganguly
South Park Mexican	http://en.wikipedia.org/wiki/South_Park_Mexican
Southern Sudan Salva Kiir	http://en.wikipedia.org/wiki/Salva_Kiir_Mayardit
Spalding Gray	http://en.wikipedia.org/wiki/Spalding_Gray
Spamford Wallace	http://en.wikipedia.org/wiki/Spamford_Wallace
Spanky McFarland	http://en.wikipedia.org/wiki/George_
Spark M. Matsunaga	http://en.wikipedia.org/wiki/Spark_M._Matsunaga
Sparky Anderson	http://en.wikipedia.org/wiki/Sparky_Anderson
Spencer Abraham	http://en.wikipedia.org/wiki/Spencer_Abraham
Spencer Bachus	http://en.wikipedia.org/wiki/Spencer_Bachus
Spencer Dryden	http://en.wikipedia.org/wiki/Spencer_Dryden
Spencer Fullerton Baird	http://en.wikipedia.org/wiki/Spencer_Fullerton_Baird
Spencer Perceval	http://en.wikipedia.org/wiki/Spencer_Perceval
Spencer Tracy	http://en.wikipedia.org/wiki/Spencer_Tracy
Spencer Tunick	http://en.wikipedia.org/wiki/Spencer_Tunick
Spice Williams	http://en.wikipedia.org/wiki/Spice_Williams
Spike Jones	http://en.wikipedia.org/wiki/Spike_Jones
Spike Jonze	http://en.wikipedia.org/wiki/Spike_Jonze
Spike Lee	http://en.wikipedia.org/wiki/Spike_Lee
Spike Milligan	http://en.wikipedia.org/wiki/Spike_Milligan
Spiro T. Agnew	http://en.wikipedia.org/wiki/Spiro_T._Agnew
Spring Byington	http://en.wikipedia.org/wiki/Spring_Byington
Squeaky Fromme	http://en.wikipedia.org/wiki/Squeaky_Fromme
Sri Chinmoy	http://en.wikipedia.org/wiki/Sri_Chinmoy
St. Agatha	http://en.wikipedia.org/wiki/St._Agatha
St. Ambrose	http://en.wikipedia.org/wiki/St._Ambrose
St. Athanasius	http://en.wikipedia.org/wiki/St._Athanasius
St. Augustine	http://en.wikipedia.org/wiki/St._Augustine
St. Augustine of Canterbury	http://en.wikipedia.org/wiki/St._Augustine_of_Canterbury
St. Bernard of Clairvaux	http://en.wikipedia.org/wiki/St._Bernard_of_Clairvaux
St. Catherine of Alexandria	http://en.wikipedia.org/wiki/St._Catherine_of_Alexandria
St. Catherine of Siena	http://en.wikipedia.org/wiki/St._Catherine_of_Siena
St. Cecilia	http://en.wikipedia.org/wiki/St._Cecilia
St. Clare	http://en.wikipedia.org/wiki/Saint_Clare_of_Assisi
St. Clement I	http://en.wikipedia.org/wiki/St._Clement_I
St. Columba	http://en.wikipedia.org/wiki/St._Columba
St. Cuthbert	http://en.wikipedia.org/wiki/St._Cuthbert
St. David	http://en.wikipedia.org/wiki/St._David
St. Denis	http://en.wikipedia.org/wiki/St._Denis
St. Dominic	http://en.wikipedia.org/wiki/St._Dominic
St. Epiphanius	http://en.wikipedia.org/wiki/Epiphanius_of_Salamis
St. Francis Borgia	http://en.wikipedia.org/wiki/St._Francis_Borgia
St. Francis de Sales	http://en.wikipedia.org/wiki/St._Francis_de_Sales
St. Francis of Assisi	http://en.wikipedia.org/wiki/St._Francis_of_Assisi
St. Francis Xavier	http://en.wikipedia.org/wiki/St._Francis_Xavier
St. George	http://en.wikipedia.org/wiki/St._George
St. Giles	http://en.wikipedia.org/wiki/St._Giles
St. Ignatius of Loyola	http://en.wikipedia.org/wiki/St._Ignatius_of_Loyola
St. Januarius	http://en.wikipedia.org/wiki/St._Januarius
St. Jerome	http://en.wikipedia.org/wiki/St._Jerome
St. John Chrysostom	http://en.wikipedia.org/wiki/St._John_Chrysostom
St. John of Beverley	http://en.wikipedia.org/wiki/John_of_Beverley
St. John of Nepomuk	http://en.wikipedia.org/wiki/St._John_of_Nepomuk
St. John of the Cross	http://en.wikipedia.org/wiki/St._John_of_the_Cross
St. Joseph	http://en.wikipedia.org/wiki/St._Joseph
St. Luke	http://en.wikipedia.org/wiki/St._Luke
St. Margaret	http://en.wikipedia.org/wiki/Saint_Margaret_of_Scotland
St. Mark	http://en.wikipedia.org/wiki/St._Mark
St. Matthew	http://en.wikipedia.org/wiki/St._Matthew
St. Nicholas	http://en.wikipedia.org/wiki/St._Nicholas
St. Oswald	http://en.wikipedia.org/wiki/Oswald_of_Northumbria
St. Peter	http://en.wikipedia.org/wiki/St._Peter
St. Philip	http://en.wikipedia.org/wiki/St._Philip
St. Pius X	http://en.wikipedia.org/wiki/St._Pius_X
St. Swithun	http://en.wikipedia.org/wiki/St._Swithun
St. Thomas Aquinas	http://en.wikipedia.org/wiki/St._Thomas_Aquinas
St. Thomas de Cantelupe	http://en.wikipedia.org/wiki/Thomas_de_Cantilupe
St. Vincent de Paul	http://en.wikipedia.org/wiki/St._Vincent_de_Paul
St. Walpurgis	http://en.wikipedia.org/wiki/Saint_Walpurga
Stacey Dash	http://en.wikipedia.org/wiki/Stacey_Dash
Stacey Grenrock-Woods	http://en.wikipedia.org/wiki/Stacey_Grenrock-Woods
Stacy Edwards	http://en.wikipedia.org/wiki/Stacy_Edwards
Stacy Ferguson	http://en.wikipedia.org/wiki/Stacy_Ferguson
Stacy Haiduk	http://en.wikipedia.org/wiki/Stacy_Haiduk
Stacy Keach	http://en.wikipedia.org/wiki/Stacy_Keach
Stan Barstow	http://en.wikipedia.org/wiki/Stan_Barstow
Stan Freberg	http://en.wikipedia.org/wiki/Stan_Freberg
Stan Getz	http://en.wikipedia.org/wiki/Stan_Getz
Stan Kenton	http://en.wikipedia.org/wiki/Stan_Kenton
Stan Laurel	http://en.wikipedia.org/wiki/Stan_Laurel
Stan Lee	http://en.wikipedia.org/wiki/Stan_Lee
Stan Lundine	http://en.wikipedia.org/wiki/Stan_Lundine
Stan Musial	http://en.wikipedia.org/wiki/Stan_Musial
Stan Parris	http://en.wikipedia.org/wiki/Stan_Parris
Stanford Moore	http://en.wikipedia.org/wiki/Stanford_Moore
Stanislao Cannizzaro	http://en.wikipedia.org/wiki/Stanislao_Cannizzaro
Stanislav Gross	http://en.wikipedia.org/wiki/Stanislav_Gross
Stanislaw Lem	http://en.wikipedia.org/wiki/Stanislaw_Lem
Stanley Baldwin	http://en.wikipedia.org/wiki/Stanley_Baldwin
Stanley Bing	http://en.wikipedia.org/wiki/Stanley_Bing
Stanley Clarke	http://en.wikipedia.org/wiki/Stanley_Clarke
Stanley Donen	http://en.wikipedia.org/wiki/Stanley_Donen
Stanley Elkin	http://en.wikipedia.org/wiki/Stanley_Elkin
Stanley Fish	http://en.wikipedia.org/wiki/Stanley_Fish
Stanley Hiller, Jr.	http://en.wikipedia.org/wiki/Stanley_Hiller
Stanley Holloway	http://en.wikipedia.org/wiki/Stanley_Holloway
Stanley Jordan	http://en.wikipedia.org/wiki/Stanley_Jordan
Stanley K. Hathaway	http://en.wikipedia.org/wiki/Stanley_K._Hathaway
Stanley Kramer	http://en.wikipedia.org/wiki/Stanley_Kramer
Stanley Kubrick	http://en.wikipedia.org/wiki/Stanley_Kubrick
Stanley Kunitz	http://en.wikipedia.org/wiki/Stanley_Kunitz
Stanley Matthews	http://en.wikipedia.org/wiki/Stanley_Matthews
Stanley Pons	http://en.wikipedia.org/wiki/Stanley_Pons
Stanley Reed	http://en.wikipedia.org/wiki/Stanley_Forman_Reed
Stanley Tucci	http://en.wikipedia.org/wiki/Stanley_Tucci
Stansfield Turner	http://en.wikipedia.org/wiki/Stansfield_Turner
Star Jones	http://en.wikipedia.org/wiki/Star_Jones
Stark Young	http://en.wikipedia.org/wiki/Stark_Young
Stedman Graham	http://en.wikipedia.org/wiki/Stedman_Graham
Steele MacKaye	http://en.wikipedia.org/wiki/Steele_MacKaye
Steen Steensen Blicher	http://en.wikipedia.org/wiki/Steen_Steensen_Blicher
Stefan George	http://en.wikipedia.org/wiki/Stefan_George
Stefanie Powers	http://en.wikipedia.org/wiki/Stefanie_Powers
Stefano Casiraghi	http://en.wikipedia.org/wiki/Stefano_Casiraghi
Stefano Della Bella	http://en.wikipedia.org/wiki/Stefano_Della_Bella
Steffi Graf	http://en.wikipedia.org/wiki/Steffi_Graf
Stella Creasy	http://en.wikipedia.org/wiki/Stella_Creasy
Stella McCartney	http://en.wikipedia.org/wiki/Stella_McCartney
Stella Stevens	http://en.wikipedia.org/wiki/Stella_Stevens
Stella Walsh	http://en.wikipedia.org/wiki/Stella_Walsh
Stellan Skarsg�rd	http://en.wikipedia.org/wiki/Stellan_Skarsg%E5rd
Sten Sture the Elder	http://en.wikipedia.org/wiki/Sten_Sture_the_Elder
Sten Sture the Younger	http://en.wikipedia.org/wiki/Sten_Sture_the_Younger
Steny H. Hoyer	http://en.wikipedia.org/wiki/Steny_H._Hoyer
Steny Hoyer	http://en.wikipedia.org/wiki/Steny_Hoyer
Stephan Brenninkmeijer	http://en.wikipedia.org/wiki/Stephan_Brenninkmeijer
Stephan Jenkins	http://en.wikipedia.org/wiki/Stephan_Jenkins
Stephan Thernstrom	http://en.wikipedia.org/wiki/Stephan_Thernstrom
St�phane Mallarm�	http://en.wikipedia.org/wiki/St%E9phane_Mallarm%E9
Stephanie Beacham	http://en.wikipedia.org/wiki/Stephanie_Beacham
Stephanie Herseth	http://en.wikipedia.org/wiki/Stephanie_Herseth
Stephanie March	http://en.wikipedia.org/wiki/Stephanie_March
Stephanie McMahon	http://en.wikipedia.org/wiki/Stephanie_McMahon
Stephanie Powers	http://en.wikipedia.org/wiki/Stephanie_Powers
Stephanie Seymour	http://en.wikipedia.org/wiki/Stephanie_Seymour
Stephanie Sun	http://en.wikipedia.org/wiki/Stephanie_Sun
Stephanie Tubbs Jones	http://en.wikipedia.org/wiki/Stephanie_Tubbs_Jones
Stephanie Zimbalist	http://en.wikipedia.org/wiki/Stephanie_Zimbalist
Stephen A. Douglas	http://en.wikipedia.org/wiki/Stephen_A._Douglas
Stephen A. Schwarzman	http://en.wikipedia.org/wiki/Stephen_A._Schwarzman
Stephen Baldwin	http://en.wikipedia.org/wiki/Stephen_Baldwin
Stephen Barclay	http://en.wikipedia.org/wiki/Stephen_Barclay
Stephen B�thory	http://en.wikipedia.org/wiki/Stephen_B%C3%A1thory_of_Poland
Stephen Blackehart	http://en.wikipedia.org/wiki/Stephen_Blackehart
Stephen Boyd	http://en.wikipedia.org/wiki/Stephen_Boyd
Stephen Breyer	http://en.wikipedia.org/wiki/Stephen_Breyer
Stephen Cambone	http://en.wikipedia.org/wiki/Stephen_Cambone
Stephen Chow	http://en.wikipedia.org/wiki/Stephen_Chow
Stephen Clark Foster	http://en.wikipedia.org/wiki/Stephen_Clark_Foster
Stephen Colbert	http://en.wikipedia.org/wiki/Stephen_Colbert
Stephen Collins	http://en.wikipedia.org/wiki/Stephen_Collins
Stephen Collins Foster	http://en.wikipedia.org/wiki/Stephen_Collins_Foster
Stephen Crabb	http://en.wikipedia.org/wiki/Stephen_Crabb
Stephen Crane	http://en.wikipedia.org/wiki/Stephen_Crane
Stephen D. Bechtel	http://en.wikipedia.org/wiki/Stephen_D._Bechtel
Stephen Decatur	http://en.wikipedia.org/wiki/Stephen_Decatur
Stephen Dorff	http://en.wikipedia.org/wiki/Stephen_Dorff
Stephen Dorrell	http://en.wikipedia.org/wiki/Stephen_Dorrell
Stephen E. Ambrose	http://en.wikipedia.org/wiki/Stephen_E._Ambrose
Stephen Fleming	http://en.wikipedia.org/wiki/Stephen_Fleming
Stephen Frears	http://en.wikipedia.org/wiki/Stephen_Frears
Stephen Fry	http://en.wikipedia.org/wiki/Stephen_Fry
Stephen Fuller Austin	http://en.wikipedia.org/wiki/Stephen_Fuller_Austin
Stephen Furst	http://en.wikipedia.org/wiki/Stephen_Furst
Stephen Gardiner	http://en.wikipedia.org/wiki/Stephen_Gardiner
Stephen Gilbert	http://en.wikipedia.org/wiki/Stephen_Gilbert_(UK_politician)
Stephen Goldsmith	http://en.wikipedia.org/wiki/Stephen_Goldsmith
Stephen Hadley	http://en.wikipedia.org/wiki/Stephen_Hadley
Stephen Hales	http://en.wikipedia.org/wiki/Stephen_Hales
Stephen Hammond	http://en.wikipedia.org/wiki/Stephen_Hammond
Stephen Harper	http://en.wikipedia.org/wiki/Stephen_Harper
Stephen Hawes	http://en.wikipedia.org/wiki/Stephen_Hawes
Stephen Hawking	http://en.wikipedia.org/wiki/Stephen_Hawking
Stephen Hepburn	http://en.wikipedia.org/wiki/Stephen_Hepburn
Stephen Hillenburg	http://en.wikipedia.org/wiki/Stephen_Hillenburg
Stephen I	http://en.wikipedia.org/wiki/Stephen_I_of_Hungary
Stephen J. Cannell	http://en.wikipedia.org/wiki/Stephen_J._Cannell
Stephen J. Solarz	http://en.wikipedia.org/wiki/Stephen_J._Solarz
Stephen Jay Gould	http://en.wikipedia.org/wiki/Stephen_Jay_Gould
Stephen King	http://en.wikipedia.org/wiki/Stephen_King
Stephen L. Neal	http://en.wikipedia.org/wiki/Stephen_L._Neal
Stephen Lang	http://en.wikipedia.org/wiki/Stephen_Lang_(actor)
Stephen Leacock	http://en.wikipedia.org/wiki/Stephen_Leacock
Stephen Lloyd	http://en.wikipedia.org/wiki/Stephen_Lloyd
Stephen Lynch	http://en.wikipedia.org/wiki/Stephen_Lynch_(politician)
Stephen M. Bennett	http://en.wikipedia.org/wiki/Steve_Bennett_(software_entrepreneur)
Stephen Malkmus	http://en.wikipedia.org/wiki/Stephen_Malkmus
Stephen Mallinder	http://en.wikipedia.org/wiki/Stephen_Mallinder
Stephen McCabe	http://en.wikipedia.org/wiki/Steve_McCabe_(politician)
Stephen McKenna	http://en.wikipedia.org/wiki/Stephen_McKenna
Stephen McPartland	http://en.wikipedia.org/wiki/Stephen_McPartland
Stephen Metcalfe	http://en.wikipedia.org/wiki/Stephen_Metcalfe_(UK_politician)
Stephen Moore	http://en.wikipedia.org/wiki/Stephen_Moore_(economist)
Stephen Moore	http://en.wikipedia.org/wiki/Stephen_Moore_(actor)
Stephen Mosley	http://en.wikipedia.org/wiki/Stephen_Mosley
Stephen Norrington	http://en.wikipedia.org/wiki/Stephen_Norrington
Stephen O'Brien	http://en.wikipedia.org/wiki/Stephen_O%27Brien
Stephen Phillips	http://en.wikipedia.org/wiki/Stephen_Phillips_(politician)
Stephen Pound	http://en.wikipedia.org/wiki/Stephen_Pound
Stephen R. Donaldson	http://en.wikipedia.org/wiki/Stephen_R._Donaldson
Stephen Rea	http://en.wikipedia.org/wiki/Stephen_Rea
Stephen Root	http://en.wikipedia.org/wiki/Stephen_Root
Stephen Solarz	http://en.wikipedia.org/wiki/Stephen_Solarz
Stephen Sommers	http://en.wikipedia.org/wiki/Stephen_Sommers
Stephen Sondheim	http://en.wikipedia.org/wiki/Stephen_Sondheim
Stephen Spender	http://en.wikipedia.org/wiki/Stephen_Spender
Stephen Stills	http://en.wikipedia.org/wiki/Stephen_Stills
Stephen Storace	http://en.wikipedia.org/wiki/Stephen_Storace
Stephen T. Early	http://en.wikipedia.org/wiki/Stephen_T._Early
Stephen Timms	http://en.wikipedia.org/wiki/Stephen_Timms
Stephen Tobolowsky	http://en.wikipedia.org/wiki/Stephen_Tobolowsky
Stephen Twigg	http://en.wikipedia.org/wiki/Stephen_Twigg
Stephen V	http://en.wikipedia.org/wiki/Stephen_V_of_Hungary
Stephen Vincent Ben�t	http://en.wikipedia.org/wiki/Stephen_Vincent_Ben%E9t
Stephen Williams	http://en.wikipedia.org/wiki/Stephen_Williams_(politician)
Stephen Wolfram	http://en.wikipedia.org/wiki/Stephen_Wolfram
Stephenson King	http://en.wikipedia.org/wiki/Stephenson_King
Stephin Merritt	http://en.wikipedia.org/wiki/Stephin_Merritt
Stepin Fetchit	http://en.wikipedia.org/wiki/Stepin_Fetchit
Sterling Hayden	http://en.wikipedia.org/wiki/Sterling_Hayden
Sterling Holloway	http://en.wikipedia.org/wiki/Sterling_Holloway
Sterling Marlin	http://en.wikipedia.org/wiki/Sterling_Marlin
Steve Albini	http://en.wikipedia.org/wiki/Steve_Albini
Steve Allen	http://en.wikipedia.org/wiki/Steve_Allen
Steve Austria	http://en.wikipedia.org/wiki/Steve_Austria
Steve Ballmer	http://en.wikipedia.org/wiki/Steve_Ballmer
Steve Barron	http://en.wikipedia.org/wiki/Steve_Barron
Steve Bartlett	http://en.wikipedia.org/wiki/Steve_Bartlett
Steve Bartman	http://en.wikipedia.org/wiki/Steve_Bartman
Steve Benen	http://en.wikipedia.org/wiki/Steve_Benen
Steve Berra	http://en.wikipedia.org/wiki/Steve_Berra
Steve Biko	http://en.wikipedia.org/wiki/Steve_Biko
Steve Bing	http://en.wikipedia.org/wiki/Steve_Bing
Steve Bloom	http://en.wikipedia.org/wiki/Steve_Bloom
Steve Brine	http://en.wikipedia.org/wiki/Steve_Brine
Steve Brodie	http://en.wikipedia.org/wiki/Steve_Brodie_(actor)
Steve Burd	http://en.wikipedia.org/wiki/Steve_Burd
Steve Burton	http://en.wikipedia.org/wiki/Steve_Burton_(actor)
Steve Buscemi	http://en.wikipedia.org/wiki/Steve_Buscemi
Steve Buyer	http://en.wikipedia.org/wiki/Steve_Buyer
Steve Carell	http://en.wikipedia.org/wiki/Steve_Carell
Steve Carlton	http://en.wikipedia.org/wiki/Steve_Carlton
Steve Case	http://en.wikipedia.org/wiki/Steve_Case
Steve Chabot	http://en.wikipedia.org/wiki/Steve_Chabot
Steve Coogan	http://en.wikipedia.org/wiki/Steve_Coogan
Steve Ditko	http://en.wikipedia.org/wiki/Steve_Ditko
Steve Driehaus	http://en.wikipedia.org/wiki/Steve_Driehaus
Steve Durand	http://en.wikipedia.org/wiki/Steve_Durand
Steve Forbes	http://en.wikipedia.org/wiki/Steve_Forbes
Steve Forrest	http://en.wikipedia.org/wiki/Steve_Forrest_(actor)
Steve Fossett	http://en.wikipedia.org/wiki/Steve_Fossett
Steve Garvey	http://en.wikipedia.org/wiki/Steve_Garvey
Steve Gibson	http://en.wikipedia.org/wiki/Steve_Gibson_(computer_programmer)
Steve Gunderson	http://en.wikipedia.org/wiki/Steve_Gunderson
Steve Guttenberg	http://en.wikipedia.org/wiki/Steve_Guttenberg
Steve Hackett	http://en.wikipedia.org/wiki/Steve_Hackett
Steve Harris	http://en.wikipedia.org/wiki/Steve_Harris_(actor)
Steve Hartman	http://en.wikipedia.org/wiki/Steve_Hartman
Steve Harvey	http://en.wikipedia.org/wiki/Steve_Harvey
Steve Hillage	http://en.wikipedia.org/wiki/Steve_Hillage
Steve Howe	http://en.wikipedia.org/wiki/Steve_Howe_(guitarist)
Steve Howe	http://en.wikipedia.org/wiki/Steve_Howe_(baseball)
Steve Irwin	http://en.wikipedia.org/wiki/Steve_Irwin
Steve Isaacs	http://en.wikipedia.org/wiki/Steve_Isaacs
Steve Israel	http://en.wikipedia.org/wiki/Steve_Israel
Steve Jackson	http://en.wikipedia.org/wiki/Steve_Jackson_(US_game_designer)
Steve Jobs	http://en.wikipedia.org/wiki/Steve_Jobs
Steve Jobs	http://en.wikipedia.org/wiki/Steve_Jobs
Steve Jones	http://en.wikipedia.org/wiki/Steve_Jones_(musician)
Steve Kagen	http://en.wikipedia.org/wiki/Steve_Kagen
Steve Kanaly	http://en.wikipedia.org/wiki/Steve_Kanaly
Steve King	http://en.wikipedia.org/wiki/Steve_King
Steve Kroft	http://en.wikipedia.org/wiki/Steve_Kroft
Steve Landesberg	http://en.wikipedia.org/wiki/Steve_Landesberg
Steve Largent	http://en.wikipedia.org/wiki/Steve_Largent
Steve Lawrence	http://en.wikipedia.org/wiki/Steve_Lawrence
Steve Lillywhite	http://en.wikipedia.org/wiki/Steve_Lillywhite
Steve Mann	http://en.wikipedia.org/wiki/Steve_Mann
Steve Mariucci	http://en.wikipedia.org/wiki/Steve_Mariucci
Steve Martin	http://en.wikipedia.org/wiki/Steve_Martin
Steve McClaren	http://en.wikipedia.org/wiki/Steve_McClaren
Steve McConnell	http://en.wikipedia.org/wiki/Steve_McConnell
Steve McQueen	http://en.wikipedia.org/wiki/Steve_McQueen
Steve Meretzky	http://en.wikipedia.org/wiki/Steve_Meretzky
Steve Miller	http://en.wikipedia.org/wiki/Steve_Miller_(musician)
Steve Miner	http://en.wikipedia.org/wiki/Steve_Miner
Steve Morse	http://en.wikipedia.org/wiki/Steve_Morse
Steve Nash	http://en.wikipedia.org/wiki/Steve_Nash
Steve Pearce	http://en.wikipedia.org/wiki/Steve_Pearce
Steve Perry	http://en.wikipedia.org/wiki/Steve_Perry_(musician)
Steve Reeves	http://en.wikipedia.org/wiki/Steve_Reeves
Steve Reich	http://en.wikipedia.org/wiki/Steve_Reich
Steve Rotheram	http://en.wikipedia.org/wiki/Steve_Rotheram
Steve Sandvoss	http://en.wikipedia.org/wiki/Steve_Sandvoss
Steve Scalise	http://en.wikipedia.org/wiki/Steve_Scalise
Steve Schiff	http://en.wikipedia.org/wiki/Steve_Schiff
Steve Swallow	http://en.wikipedia.org/wiki/Steve_Swallow
Steve Symms	http://en.wikipedia.org/wiki/Steve_Symms
Steve Vai	http://en.wikipedia.org/wiki/Steve_Vai
Steve Van Zandt	http://en.wikipedia.org/wiki/Steve_Van_Zandt
Steve Watson	http://en.wikipedia.org/wiki/Steve_Watson_(actor)
Steve Webb	http://en.wikipedia.org/wiki/Steve_Webb
Steve Winwood	http://en.wikipedia.org/wiki/Steve_Winwood
Steve Wozniak	http://en.wikipedia.org/wiki/Steve_Wozniak
Steve Wynn	http://en.wikipedia.org/wiki/Steve_Wynn_(entrepreneur)
Steve Young	http://en.wikipedia.org/wiki/Steve_Young_(American_football)
Steve Zahn	http://en.wikipedia.org/wiki/Steve_Zahn
Steven A. Ballmer	http://en.wikipedia.org/wiki/Steven_A._Ballmer
Steven A. Burd	http://en.wikipedia.org/wiki/Steven_Burd
Steven Adler	http://en.wikipedia.org/wiki/Steven_Adler
Steven Baker	http://en.wikipedia.org/wiki/Steve_Baker_(UK_politician)
Steven Bauer	http://en.wikipedia.org/wiki/Steven_Bauer
Steven Berkoff	http://en.wikipedia.org/wiki/Steven_Berkoff
Steven Bochco	http://en.wikipedia.org/wiki/Steven_Bochco
Steven Chu	http://en.wikipedia.org/wiki/Steven_Chu
Steven Cojocaru	http://en.wikipedia.org/wiki/Steven_Cojocaru
Steven Culp	http://en.wikipedia.org/wiki/Steven_Culp
Steven Drozd	http://en.wikipedia.org/wiki/Steven_Drozd
Steven Gerrard	http://en.wikipedia.org/wiki/Steven_Gerrard
Steven Hatfill	http://en.wikipedia.org/wiki/Steven_Hatfill
Steven Hill	http://en.wikipedia.org/wiki/Steven_Hill
Steven Hoefflin	http://en.wikipedia.org/wiki/Steven_Hoefflin
Steven Jesse Bernstein	http://en.wikipedia.org/wiki/Steven_Jesse_Bernstein
Steven LaTourette	http://en.wikipedia.org/wiki/Steven_LaTourette
Steven Levitt	http://en.wikipedia.org/wiki/Steven_Levitt
Steven Levy	http://en.wikipedia.org/wiki/Steven_Levy
Steven M. Bornstein	http://en.wikipedia.org/wiki/Steve_Bornstein
Steven Michaels	http://en.wikipedia.org/wiki/Steven_Michaels
Steven Millhauser	http://en.wikipedia.org/wiki/Steven_Millhauser
Steven Pinker	http://en.wikipedia.org/wiki/Steven_Pinker
Steven Rothman	http://en.wikipedia.org/wiki/Steven_Rothman
Steven Seagal	http://en.wikipedia.org/wiki/Steven_Seagal
Steven Soderbergh	http://en.wikipedia.org/wiki/Steven_Soderbergh
Steven Spielberg	http://en.wikipedia.org/wiki/Steven_Spielberg
Steven Stapleton	http://en.wikipedia.org/wiki/Steven_Stapleton
Steven Stayner	http://en.wikipedia.org/wiki/Steven_Stayner
Steven T. Katz	http://en.wikipedia.org/wiki/Steven_T._Katz
Steven Tyler	http://en.wikipedia.org/wiki/Steven_Tyler
Steven Weber	http://en.wikipedia.org/wiki/Steven_Weber_(actor)
Steven Weinberg	http://en.wikipedia.org/wiki/Steven_Weinberg
Steven Wright	http://en.wikipedia.org/wiki/Steven_Wright
Stevie Nicks	http://en.wikipedia.org/wiki/Stevie_Nicks
Stevie Ray Vaughan	http://en.wikipedia.org/wiki/Stevie_Ray_Vaughan
Stevie Wonder	http://en.wikipedia.org/wiki/Stevie_Wonder
Stew Albert	http://en.wikipedia.org/wiki/Stew_Albert
Stewart B. McKinney	http://en.wikipedia.org/wiki/Stewart_B._McKinney
Stewart Brand	http://en.wikipedia.org/wiki/Stewart_Brand
Stewart Copeland	http://en.wikipedia.org/wiki/Stewart_Copeland
Stewart Granger	http://en.wikipedia.org/wiki/Stewart_Granger
Stewart Hosie	http://en.wikipedia.org/wiki/Stewart_Hosie
Stewart Jackson	http://en.wikipedia.org/wiki/Stewart_Jackson
Stewart Udall	http://en.wikipedia.org/wiki/Stewart_Udall
Sticky Fingaz	http://en.wikipedia.org/wiki/Sticky_Fingaz
Stjepan Mesic	http://en.wikipedia.org/wiki/Stjepan_Mesic
Stjepan Mesic	http://en.wikipedia.org/wiki/Stjepan_Mesic
Stockard Channing	http://en.wikipedia.org/wiki/Stockard_Channing
Stokely Carmichael	http://en.wikipedia.org/wiki/Stokely_Carmichael
Stone Cold Steve Austin	http://en.wikipedia.org/wiki/Stone_Cold_Steve_Austin
Stone Gossard	http://en.wikipedia.org/wiki/Stone_Gossard
Stone Phillips	http://en.wikipedia.org/wiki/Stone_Phillips
Stonewall Jackson	http://en.wikipedia.org/wiki/Stonewall_Jackson
Storm Jameson	http://en.wikipedia.org/wiki/Storm_Jameson
Story Musgrave	http://en.wikipedia.org/wiki/Story_Musgrave
Strobe Talbott	http://en.wikipedia.org/wiki/Strobe_Talbott
Strom Thurmond	http://en.wikipedia.org/wiki/Strom_Thurmond
Strom Thurmond	http://en.wikipedia.org/wiki/Strom_Thurmond
Strother Martin	http://en.wikipedia.org/wiki/Strother_Martin
Stu Phillips	http://en.wikipedia.org/wiki/Stu_Phillips_(composer)
Stuart Adamson	http://en.wikipedia.org/wiki/Stuart_Adamson
Stuart Andrew	http://en.wikipedia.org/wiki/Stuart_Andrew
Stuart Bell	http://en.wikipedia.org/wiki/Stuart_Bell
Stuart Davis	http://en.wikipedia.org/wiki/Stuart_Davis_(painter)
Stuart Elliott	http://en.wikipedia.org/wiki/Stuart_Elliott_(drummer)
Stuart Margolin	http://en.wikipedia.org/wiki/Stuart_Margolin
Stuart Murdoch	http://en.wikipedia.org/wiki/Stuart_Murdoch_(musician)
Stuart Rosenberg	http://en.wikipedia.org/wiki/Stuart_Rosenberg
Stuart Sutcliffe	http://en.wikipedia.org/wiki/Stuart_Sutcliffe
Stuart Symington	http://en.wikipedia.org/wiki/Stuart_Symington
Stuart Townsend	http://en.wikipedia.org/wiki/Stuart_Townsend
Stuart Whitman	http://en.wikipedia.org/wiki/Stuart_Whitman
Stubby Kaye	http://en.wikipedia.org/wiki/Stubby_Kaye
Studs Terkel	http://en.wikipedia.org/wiki/Studs_Terkel
Stuttering John	http://en.wikipedia.org/wiki/Stuttering_John
Su Tseng-chang	http://en.wikipedia.org/wiki/Su_Tseng-chang
Subcomandante Marcos	http://en.wikipedia.org/wiki/Subcomandante_Marcos
Subrahmanyan Chandrasekhar	http://en.wikipedia.org/wiki/Subrahmanyan_Chandrasekhar
Sue Grafton	http://en.wikipedia.org/wiki/Sue_Grafton
Sue Johanson	http://en.wikipedia.org/wiki/Sue_Johanson
Sue Kelly	http://en.wikipedia.org/wiki/Sue_Kelly
Sue Lyon	http://en.wikipedia.org/wiki/Sue_Lyon
Sue Myrick	http://en.wikipedia.org/wiki/Sue_Myrick
Suehiro Maruo	http://en.wikipedia.org/wiki/Suehiro_Maruo
Sugar Ray Leonard	http://en.wikipedia.org/wiki/Sugar_Ray_Leonard
Sugar Ray Robinson	http://en.wikipedia.org/wiki/Sugar_Ray_Robinson
Suge Knight	http://en.wikipedia.org/wiki/Suge_Knight
S�khbaataryn Batbold	http://en.wikipedia.org/wiki/S%FCkhbaataryn_Batbold
Suleiman II	http://en.wikipedia.org/wiki/Suleiman_II
Suleiman the Magnificent	http://en.wikipedia.org/wiki/Suleiman_the_Magnificent
Sully Erna	http://en.wikipedia.org/wiki/Sully_Erna
Sully Prudhomme	http://en.wikipedia.org/wiki/Sully_Prudhomme
Summer Phoenix	http://en.wikipedia.org/wiki/Summer_Phoenix
Summer Sanders	http://en.wikipedia.org/wiki/Summer_Sanders
Sumner Redstone	http://en.wikipedia.org/wiki/Sumner_Redstone
Sun Myung Moon	http://en.wikipedia.org/wiki/Sun_Myung_Moon
Sun Ra	http://en.wikipedia.org/wiki/Sun_Ra
Sun Tzu	http://en.wikipedia.org/wiki/Sun_Tzu
Sun Yat-sen	http://en.wikipedia.org/wiki/Sun_Yat-sen
Sunil Gavaskar	http://en.wikipedia.org/wiki/Sunil_Gavaskar
Sunny Deol	http://en.wikipedia.org/wiki/Sunny_Deol
Sunny Murray	http://en.wikipedia.org/wiki/Sunny_Murray
Sunny von Bulow	http://en.wikipedia.org/wiki/Sunny_von_Bulow
Super Cat	http://en.wikipedia.org/wiki/Super_Cat
Super Dave Osborne	http://en.wikipedia.org/wiki/Super_Dave_Osborne
Suraj ud Dowlah	http://en.wikipedia.org/wiki/Siraj_ud-Daulah
Susan Anspach	http://en.wikipedia.org/wiki/Susan_Anspach
Susan Anton	http://en.wikipedia.org/wiki/Susan_Anton
Susan B. Anthony	http://en.wikipedia.org/wiki/Susan_B._Anthony
Susan Blackmore	http://en.wikipedia.org/wiki/Susan_Blackmore
Susan Blakely	http://en.wikipedia.org/wiki/Susan_Blakely
Susan Block	http://en.wikipedia.org/wiki/Susan_Block
Susan Collins	http://en.wikipedia.org/wiki/Susan_Collins
Susan Coolidge	http://en.wikipedia.org/wiki/Susan_Coolidge
Susan Davis	http://en.wikipedia.org/wiki/Susan_Davis_(Congresswoman)
Susan Dey	http://en.wikipedia.org/wiki/Susan_Dey
Susan Estrich	http://en.wikipedia.org/wiki/Susan_Estrich
Susan Faludi	http://en.wikipedia.org/wiki/Susan_Faludi
Susan Flannery	http://en.wikipedia.org/wiki/Susan_Flannery
Susan George	http://en.wikipedia.org/wiki/Susan_George_(actress)
Susan Glaspell	http://en.wikipedia.org/wiki/Susan_Glaspell
Susan Hampshire	http://en.wikipedia.org/wiki/Susan_Hampshire
Susan Hayward	http://en.wikipedia.org/wiki/Susan_Hayward
Susan Jacoby	http://en.wikipedia.org/wiki/Susan_Jacoby
Susan Jones	http://en.wikipedia.org/wiki/Susan_Jones
Susan Lucci	http://en.wikipedia.org/wiki/Susan_Lucci
Susan McDougal	http://en.wikipedia.org/wiki/Susan_McDougal
Susan Oliver	http://en.wikipedia.org/wiki/Susan_Oliver
Susan Olsen	http://en.wikipedia.org/wiki/Susan_Olsen
Susan Powter	http://en.wikipedia.org/wiki/Susan_Powter
Susan Saint James	http://en.wikipedia.org/wiki/Susan_Saint_James
Susan Sarandon	http://en.wikipedia.org/wiki/Susan_Sarandon
Susan Sontag	http://en.wikipedia.org/wiki/Susan_Sontag
Susan St. James	http://en.wikipedia.org/wiki/Susan_St._James
Susan Sullivan	http://en.wikipedia.org/wiki/Susan_Sullivan
Susan Tyrrell	http://en.wikipedia.org/wiki/Susan_Tyrrell
Susan Ward	http://en.wikipedia.org/wiki/Susan_Ward
Susanna Hoffs	http://en.wikipedia.org/wiki/Susanna_Hoffs
Susanna Rowson	http://en.wikipedia.org/wiki/Susanna_Rowson
Susanne Alfvengren	http://en.wikipedia.org/wiki/Susanne_Alfvengren
Susie Bright	http://en.wikipedia.org/wiki/Susie_Bright
Susilo Bambang Yudhoyono	http://en.wikipedia.org/wiki/Susilo_Bambang_Yudhoyono
Suzanne Kosmas	http://en.wikipedia.org/wiki/Suzanne_Kosmas
Suzanne Pleshette	http://en.wikipedia.org/wiki/Suzanne_Pleshette
Suzanne Somers	http://en.wikipedia.org/wiki/Suzanne_Somers
Suzanne Vega	http://en.wikipedia.org/wiki/Suzanne_Vega
Suze Orman	http://en.wikipedia.org/wiki/Suze_Orman
Suze Randall	http://en.wikipedia.org/wiki/Suze_Randall
Suzi Quatro	http://en.wikipedia.org/wiki/Suzi_Quatro
Suzy Aiken	http://en.wikipedia.org/wiki/Suzy_Aiken
Suzy Amis	http://en.wikipedia.org/wiki/Suzy_Amis
Suzy Chaffee	http://en.wikipedia.org/wiki/Suzy_Chaffee
Svante Arrhenius	http://en.wikipedia.org/wiki/Svante_Arrhenius
Sven-Goran Eriksson	http://en.wikipedia.org/wiki/Sven-Goran_Eriksson
Svetozar Marovic	http://en.wikipedia.org/wiki/Svetozar_Marovic
Sweetie Irie	http://en.wikipedia.org/wiki/Sweetie_Irie
Sweyn Forkbeard	http://en.wikipedia.org/wiki/Sweyn_Forkbeard
Swoosie Kurtz	http://en.wikipedia.org/wiki/Swoosie_Kurtz
Sybille Bedford	http://en.wikipedia.org/wiki/Sybille_Bedford
Syd Barrett	http://en.wikipedia.org/wiki/Syd_Barrett
Syd Hoff	http://en.wikipedia.org/wiki/Syd_Hoff
Syd Straw	http://en.wikipedia.org/wiki/Syd_Straw
Sydney Greenstreet	http://en.wikipedia.org/wiki/Sydney_Greenstreet
Sydney Penny	http://en.wikipedia.org/wiki/Sydney_Penny
Sydney Pollack	http://en.wikipedia.org/wiki/Sydney_Pollack
Sydney Schanberg	http://en.wikipedia.org/wiki/Sydney_Schanberg
Sydney Smith	http://en.wikipedia.org/wiki/Sydney_Smith
Sylvester Stallone	http://en.wikipedia.org/wiki/Sylvester_Stallone
Sylvia Ashton-Warner	http://en.wikipedia.org/wiki/Sylvia_Ashton-Warner
Sylvia Browne	http://en.wikipedia.org/wiki/Sylvia_Browne
Sylvia Hermon	http://en.wikipedia.org/wiki/Sylvia_Hermon
Sylvia Plath	http://en.wikipedia.org/wiki/Sylvia_Plath
Sylvia Sidney	http://en.wikipedia.org/wiki/Sylvia_Sidney
Sylvia Syms	http://en.wikipedia.org/wiki/Sylvia_Syms
Sylvia Townsend Warner	http://en.wikipedia.org/wiki/Sylvia_Townsend_Warner
Symeon Metaphrastes	http://en.wikipedia.org/wiki/Symeon_Metaphrastes
Syngman Rhee	http://en.wikipedia.org/wiki/Syngman_Rhee
Szolem Mandelbrojt	http://en.wikipedia.org/wiki/Szolem_Mandelbrojt
T. Boone Pickens	http://en.wikipedia.org/wiki/T._Boone_Pickens
T. C. Boyle	http://en.wikipedia.org/wiki/T._C._Boyle
T. D. Jakes	http://en.wikipedia.org/wiki/T._D._Jakes
T. E. Lawrence	http://en.wikipedia.org/wiki/T._E._Lawrence
T. H. White	http://en.wikipedia.org/wiki/T._H._White
T. I.	http://en.wikipedia.org/wiki/T._I.
T. M. Aluko	http://en.wikipedia.org/wiki/T._M._Aluko
T. S. Eliot	http://en.wikipedia.org/wiki/T._S._Eliot
T. S. Stribling	http://en.wikipedia.org/wiki/T._S._Stribling
Tab Hunter	http://en.wikipedia.org/wiki/Tab_Hunter
Tabar� Ram�n V�zquez Rosas	http://en.wikipedia.org/wiki/Tabar%E9_Ram%F3n_V%E1zquez_Rosas
Tabitha Soren	http://en.wikipedia.org/wiki/Tabitha_Soren
Tadeusz Borowski	http://en.wikipedia.org/wiki/Tadeusz_Borowski
Tadeusz Kosciuszko	http://en.wikipedia.org/wiki/Tadeusz_Kosciuszko
Taher Elgamal	http://en.wikipedia.org/wiki/Taher_Elgamal
Tahj Mowry	http://en.wikipedia.org/wiki/Tahj_Mowry
Tahnee Welch	http://en.wikipedia.org/wiki/Tahnee_Welch
Tai Babilonia	http://en.wikipedia.org/wiki/Tai_Babilonia
Taisuke Itagaki	http://en.wikipedia.org/wiki/Taisuke_Itagaki
Takashi Miike	http://en.wikipedia.org/wiki/Takashi_Miike
Takeuchi Naoko	http://en.wikipedia.org/wiki/Takeuchi_Naoko
Talcott Parsons	http://en.wikipedia.org/wiki/Talcott_Parsons
Talia Shire	http://en.wikipedia.org/wiki/Talia_Shire
Talib Kweli	http://en.wikipedia.org/wiki/Talib_Kweli
Talisa Soto	http://en.wikipedia.org/wiki/Talisa_Soto
Tallulah Bankhead	http://en.wikipedia.org/wiki/Tallulah_Bankhead
Talvin Singh	http://en.wikipedia.org/wiki/Talvin_Singh
Talwinder Singh Parmar	http://en.wikipedia.org/wiki/Talwinder_Singh_Parmar
Tam White	http://en.wikipedia.org/wiki/Tam_White
Tamera Mowry	http://en.wikipedia.org/wiki/Tamera_Mowry
Tammi Terrell	http://en.wikipedia.org/wiki/Tammi_Terrell
Tammy Baldwin	http://en.wikipedia.org/wiki/Tammy_Baldwin
Tammy Blanchard	http://en.wikipedia.org/wiki/Tammy_Blanchard
Tammy Bruce	http://en.wikipedia.org/wiki/Tammy_Bruce
Tammy Duckworth	http://en.wikipedia.org/wiki/Tammy_Duckworth
Tammy Faye Bakker	http://en.wikipedia.org/wiki/Tammy_Faye_Bakker
Tammy Grimes	http://en.wikipedia.org/wiki/Tammy_Grimes
Tammy Lynn Michaels	http://en.wikipedia.org/wiki/Tammy_Lynn_Michaels
Tammy Wynette	http://en.wikipedia.org/wiki/Tammy_Wynette
Tandja Mamadou	http://en.wikipedia.org/wiki/Tandja_Mamadou
Tantia Topi	http://en.wikipedia.org/wiki/Tantia_Topi
Tanya Allen	http://en.wikipedia.org/wiki/Tanya_Allen
Tanya Donelly	http://en.wikipedia.org/wiki/Tanya_Donelly
Tanya Roberts	http://en.wikipedia.org/wiki/Tanya_Roberts
Tanya Tagaq Gillis	http://en.wikipedia.org/wiki/Tanya_Tagaq_Gillis
Tanya Tucker	http://en.wikipedia.org/wiki/Tanya_Tucker
Tara Lipinski	http://en.wikipedia.org/wiki/Tara_Lipinski
Tara Reid	http://en.wikipedia.org/wiki/Tara_Reid
Tara Strong	http://en.wikipedia.org/wiki/Tara_Strong
Taran Noah Smith	http://en.wikipedia.org/wiki/Taran_Noah_Smith
Tariq al-Hashimi	http://en.wikipedia.org/wiki/Tariq_al-Hashimi
Tariq Aziz	http://en.wikipedia.org/wiki/Tariq_Aziz
Tarja Halonen	http://en.wikipedia.org/wiki/Tarja_Halonen
Tarquinius Priscus	http://en.wikipedia.org/wiki/Tarquinius_Priscus
Tarquinius Superbus	http://en.wikipedia.org/wiki/Tarquinius_Superbus
Taryn Manning	http://en.wikipedia.org/wiki/Taryn_Manning
Tassos Papadopoulos	http://en.wikipedia.org/wiki/Tassos_Papadopoulos
Tate Donovan	http://en.wikipedia.org/wiki/Tate_Donovan
Tatjana Patitz	http://en.wikipedia.org/wiki/Tatjana_Patitz
Tatum O'Neal	http://en.wikipedia.org/wiki/Tatum_O%27Neal
Tatyana Ali	http://en.wikipedia.org/wiki/Tatyana_Ali
Taufa'ahau Tupou IV	http://en.wikipedia.org/wiki/Taufa%27ahau_Tupou_IV
Tavis Smiley	http://en.wikipedia.org/wiki/Tavis_Smiley
Tawny Kitaen	http://en.wikipedia.org/wiki/Tawny_Kitaen
Tay Garnett	http://en.wikipedia.org/wiki/Tay_Garnett
Taye Diggs	http://en.wikipedia.org/wiki/Taye_Diggs
Taylor Dayne	http://en.wikipedia.org/wiki/Taylor_Dayne
Taylor Hackford	http://en.wikipedia.org/wiki/Taylor_Hackford
Taylor Hanson	http://en.wikipedia.org/wiki/Taylor_Hanson
Taylor Hawkins	http://en.wikipedia.org/wiki/Taylor_Hawkins
Taylor Negron	http://en.wikipedia.org/wiki/Taylor_Negron
T-Bone Burnett	http://en.wikipedia.org/wiki/T-Bone_Burnett
T-Bone Walker	http://en.wikipedia.org/wiki/T-Bone_Walker
Tea Leoni	http://en.wikipedia.org/wiki/Tea_Leoni
Tea Leoni	http://en.wikipedia.org/wiki/Tea_Leoni
Ted Allen	http://en.wikipedia.org/wiki/Ted_Allen
Ted Allen	http://en.wikipedia.org/wiki/Ted_Allen
Ted Bessell	http://en.wikipedia.org/wiki/Ted_Bessell
Ted Bundy	http://en.wikipedia.org/wiki/Ted_Bundy
Ted Cassidy	http://en.wikipedia.org/wiki/Ted_Cassidy
Ted Danson	http://en.wikipedia.org/wiki/Ted_Danson
Ted Demme	http://en.wikipedia.org/wiki/Ted_Demme
Ted Deutch	http://en.wikipedia.org/wiki/Ted_Deutch
Ted Hughes	http://en.wikipedia.org/wiki/Ted_Hughes
Ted Kaczynski	http://en.wikipedia.org/wiki/Ted_Kaczynski
Ted Kaufman	http://en.wikipedia.org/wiki/Ted_Kaufman
Ted Kennedy	http://en.wikipedia.org/wiki/Ted_Kennedy
Ted Knight	http://en.wikipedia.org/wiki/Ted_Knight
Ted Kooser	http://en.wikipedia.org/wiki/Ted_Kooser
Ted Koppel	http://en.wikipedia.org/wiki/Ted_Koppel
Ted Kotcheff	http://en.wikipedia.org/wiki/Ted_Kotcheff
Ted Kulongoski	http://en.wikipedia.org/wiki/Ted_Kulongoski
Ted Lange	http://en.wikipedia.org/wiki/Ted_Lange
Ted Levine	http://en.wikipedia.org/wiki/Ted_Levine
Ted Lindsay	http://en.wikipedia.org/wiki/Ted_Lindsay
Ted McGinley	http://en.wikipedia.org/wiki/Ted_McGinley
Ted Nelson	http://en.wikipedia.org/wiki/Ted_Nelson
Ted Nugent	http://en.wikipedia.org/wiki/Ted_Nugent
Ted Olson	http://en.wikipedia.org/wiki/Theodore_Olson
Ted Poe	http://en.wikipedia.org/wiki/Ted_Poe
Ted Radcliffe	http://en.wikipedia.org/wiki/Ted_Radcliffe
Ted Rall	http://en.wikipedia.org/wiki/Ted_Rall
Ted Ross	http://en.wikipedia.org/wiki/Ted_Ross
Ted Schroeder	http://en.wikipedia.org/wiki/Ted_Schroeder
Ted Sorensen	http://en.wikipedia.org/wiki/Ted_Sorensen
Ted Stevens	http://en.wikipedia.org/wiki/Ted_Stevens
Ted Strickland	http://en.wikipedia.org/wiki/Ted_Strickland
Ted Turner	http://en.wikipedia.org/wiki/Ted_Turner
Ted Wass	http://en.wikipedia.org/wiki/Ted_Wass_(actor)
Ted Weiss	http://en.wikipedia.org/wiki/Ted_Weiss
Ted Williams	http://en.wikipedia.org/wiki/Ted_Williams
Teddy Pendergrass	http://en.wikipedia.org/wiki/Teddy_Pendergrass
Teddy Riley	http://en.wikipedia.org/wiki/Teddy_Riley_(producer)
Teemu Aalto	http://en.wikipedia.org/wiki/Teemu_Aalto
Teena Marie	http://en.wikipedia.org/wiki/Teena_Marie
Tego Calder�n	http://en.wikipedia.org/wiki/Tego_Calder%F3n
Telly Savalas	http://en.wikipedia.org/wiki/Telly_Savalas
Telma Hopkins	http://en.wikipedia.org/wiki/Telma_Hopkins
Tempestt Bledsoe	http://en.wikipedia.org/wiki/Tempestt_Bledsoe
Temple Grandin	http://en.wikipedia.org/wiki/Temple_Grandin
Tengai Amano	http://en.wikipedia.org/wiki/Tengai_Amano
Tennessee Ernie Ford	http://en.wikipedia.org/wiki/Tennessee_Ernie_Ford
Tennessee Williams	http://en.wikipedia.org/wiki/Tennessee_Williams
Tenzing Norgay	http://en.wikipedia.org/wiki/Tenzing_Norgay
Teodoro Obiang Nguema Mbasogo	http://en.wikipedia.org/wiki/Teodoro_Obiang_Nguema_Mbasogo
Terence Fisher	http://en.wikipedia.org/wiki/Terence_Fisher
Terence Hill	http://en.wikipedia.org/wiki/Terence_Hill
Terence McKenna	http://en.wikipedia.org/wiki/Terence_McKenna
Terence Rattigan	http://en.wikipedia.org/wiki/Terence_Rattigan
Terence Stamp	http://en.wikipedia.org/wiki/Terence_Stamp
Terence Trent D'Arby	http://en.wikipedia.org/wiki/Terence_Trent_D%27Arby
Terence Young	http://en.wikipedia.org/wiki/Terence_Young_(director)
Teresa Heinz	http://en.wikipedia.org/wiki/Teresa_Heinz
Teresa Pearce	http://en.wikipedia.org/wiki/Teresa_Pearce
Teresa Wright	http://en.wikipedia.org/wiki/Teresa_Wright
Teri Garr	http://en.wikipedia.org/wiki/Teri_Garr
Teri Hatcher	http://en.wikipedia.org/wiki/Teri_Hatcher
Teri Polo	http://en.wikipedia.org/wiki/Teri_Polo
Terrance Stamp	http://en.wikipedia.org/wiki/Terrance_Stamp
Terrell Owens	http://en.wikipedia.org/wiki/Terrell_Owens
Terrence Howard	http://en.wikipedia.org/wiki/Terrence_Howard
Terrence Malick	http://en.wikipedia.org/wiki/Terrence_Malick
Terrence McNally	http://en.wikipedia.org/wiki/Terrence_McNally
Terri Clark	http://en.wikipedia.org/wiki/Terri_Clark
Terri Schiavo	http://en.wikipedia.org/wiki/Terri_Schiavo
Terry Allen	http://en.wikipedia.org/wiki/Terry_Allen_%28American_football_coach%29
Terry Bozzio	http://en.wikipedia.org/wiki/Terry_Bozzio
Terry Bradshaw	http://en.wikipedia.org/wiki/Terry_Bradshaw
Terry Brooks	http://en.wikipedia.org/wiki/Terry_Brooks
Terry Crews	http://en.wikipedia.org/wiki/Terry_Crews
Terry Everett	http://en.wikipedia.org/wiki/Terry_Everett
Terry Farrell	http://en.wikipedia.org/wiki/Terry_Farrell_(actress)
Terry Gilliam	http://en.wikipedia.org/wiki/Terry_Gilliam
Terry Goodkind	http://en.wikipedia.org/wiki/Terry_Goodkind
Terry Gross	http://en.wikipedia.org/wiki/Terry_Gross
Terry J. Lundgren	http://en.wikipedia.org/wiki/Terry_J._Lundgren
Terry Jones	http://en.wikipedia.org/wiki/Terry_Jones
Terry L. Bruce	http://en.wikipedia.org/wiki/Terry_L._Bruce
Terry Lanni	http://en.wikipedia.org/wiki/Terrence_Lanni
Terry McAuliffe	http://en.wikipedia.org/wiki/Terry_McAuliffe
Terry McGuirk	http://en.wikipedia.org/wiki/Terry_McGuirk
Terry McMillan	http://en.wikipedia.org/wiki/Terry_McMillan
Terry Melcher	http://en.wikipedia.org/wiki/Terry_Melcher
Terry Moore	http://en.wikipedia.org/wiki/Terry_Moore_(actress)
Terry Moran	http://en.wikipedia.org/wiki/Terry_Moran
Terry Nichols	http://en.wikipedia.org/wiki/Terry_Nichols
Terry O'Quinn	http://en.wikipedia.org/wiki/Terry_O%27Quinn
Terry Pratchett	http://en.wikipedia.org/wiki/Terry_Pratchett
Terry Riley	http://en.wikipedia.org/wiki/Terry_Riley
Terry Sanford	http://en.wikipedia.org/wiki/Terry_Sanford
Terry Semel	http://en.wikipedia.org/wiki/Terry_Semel
Terry Waite	http://en.wikipedia.org/wiki/Terry_Waite
Terry Winograd	http://en.wikipedia.org/wiki/Terry_Winograd
Terry Wogan	http://en.wikipedia.org/wiki/Terry_Wogan
Terry Zwigoff	http://en.wikipedia.org/wiki/Terry_Zwigoff
Tertius Zongo	http://en.wikipedia.org/wiki/Tertius_Zongo
Tessa Allen	http://en.wikipedia.org/wiki/Tessa_Allen
Tessa Jowell	http://en.wikipedia.org/wiki/Tessa_Jowell
Tessa Munt	http://en.wikipedia.org/wiki/Tessa_Munt
Tetsuro Amino	http://en.wikipedia.org/wiki/Tetsuro_Amino
Tevin Campbell	http://en.wikipedia.org/wiki/Tevin_Campbell
Tewfik Pasha	http://en.wikipedia.org/wiki/Tewfik_Pasha
Tex Avery	http://en.wikipedia.org/wiki/Tex_Avery
Tex Ritter	http://en.wikipedia.org/wiki/Tex_Ritter
Tex Schramm	http://en.wikipedia.org/wiki/Tex_Schramm
Tex Watson	http://en.wikipedia.org/wiki/Tex_Watson
Thabo Mbeki	http://en.wikipedia.org/wiki/Thabo_Mbeki
Thabo Mbeki	http://en.wikipedia.org/wiki/Thabo_Mbeki
Thad Allen	http://en.wikipedia.org/wiki/Thad_Allen
Thad Cochran	http://en.wikipedia.org/wiki/Thad_Cochran
Thad Cochran	http://en.wikipedia.org/wiki/Thad_Cochran
Thad Jones	http://en.wikipedia.org/wiki/Thad_Jones
Thaddeus McCotter	http://en.wikipedia.org/wiki/Thaddeus_McCotter
Thaddeus Stevens	http://en.wikipedia.org/wiki/Thaddeus_Stevens
Thaksin Shinawatra	http://en.wikipedia.org/wiki/Thaksin_Shinawatra
Than Shwe	http://en.wikipedia.org/wiki/Than_Shwe
Than Shwe	http://en.wikipedia.org/wiki/Than_Shwe
Thandie Newton	http://en.wikipedia.org/wiki/Thandie_Newton
Thayer David	http://en.wikipedia.org/wiki/Thayer_David
The B�b	http://en.wikipedia.org/wiki/The_B%E1b
The Legendary Stardust Cowboy	http://en.wikipedia.org/wiki/The_Legendary_Stardust_Cowboy
The Madd Rapper	http://en.wikipedia.org/wiki/The_Madd_Rapper
The Michael Toy	http://en.wikipedia.org/wiki/Michael_Toy
The RZA	http://en.wikipedia.org/wiki/The_RZA
The Svedberg	http://en.wikipedia.org/wiki/The_Svedberg
Thea Astley	http://en.wikipedia.org/wiki/Thea_Astley
Thea Gill	http://en.wikipedia.org/wiki/Thea_Gill
Theda Bara	http://en.wikipedia.org/wiki/Theda_Bara
Thein Sein	http://en.wikipedia.org/wiki/Thein_Sein
Thelma Drake	http://en.wikipedia.org/wiki/Thelma_Drake
Thelma Ritter	http://en.wikipedia.org/wiki/Thelma_Ritter
Thelma Todd	http://en.wikipedia.org/wiki/Thelma_Todd
Thelonious Monk	http://en.wikipedia.org/wiki/Thelonious_Monk
Themba Dlamini	http://en.wikipedia.org/wiki/Themba_Dlamini
Theo Albrecht	http://en.wikipedia.org/wiki/Theo_Albrecht
Theo de Raadt	http://en.wikipedia.org/wiki/Theo_de_Raadt
Theo Epstein	http://en.wikipedia.org/wiki/Theo_Epstein
Theo Van Gogh	http://en.wikipedia.org/wiki/Theo_van_Gogh_(film_director)
Theobald von Bethmann-Hollweg	http://en.wikipedia.org/wiki/Theobald_von_Bethmann-Hollweg
Theodor Adorno	http://en.wikipedia.org/wiki/Theodor_Adorno
Theodor Billroth	http://en.wikipedia.org/wiki/Theodor_Billroth
Theodor de Bry	http://en.wikipedia.org/wiki/Theodor_de_Bry
Theodor Fontane	http://en.wikipedia.org/wiki/Theodor_Fontane
Theodor Herzl	http://en.wikipedia.org/wiki/Theodor_Herzl
Theodor Heuss	http://en.wikipedia.org/wiki/Theodor_Heuss
Theodor Mommsen	http://en.wikipedia.org/wiki/Theodor_Mommsen
Theodor Reuss	http://en.wikipedia.org/wiki/Theodor_Reuss
Theodor Schwann	http://en.wikipedia.org/wiki/Theodor_Schwann
Theodor Storm	http://en.wikipedia.org/wiki/Theodor_Storm
Theodore Beza	http://en.wikipedia.org/wiki/Theodore_Beza
Theodore Bikel	http://en.wikipedia.org/wiki/Theodore_Bikel
Theodore Dreiser	http://en.wikipedia.org/wiki/Theodore_Dreiser
Theodore F. Stevens	http://en.wikipedia.org/wiki/Theodore_F._Stevens
Th�odore G�ricault	http://en.wikipedia.org/wiki/Th%E9odore_G%E9ricault
Theodore H. White	http://en.wikipedia.org/wiki/Theodore_H._White
Theodore Roethke	http://en.wikipedia.org/wiki/Theodore_Roethke
Theodore Roosevelt	http://en.wikipedia.org/wiki/Theodore_Roosevelt
Th�odore Rousseau	http://en.wikipedia.org/wiki/Th%E9odore_Rousseau
Theodore Sturgeon	http://en.wikipedia.org/wiki/Theodore_Sturgeon
Theodore W. Richards	http://en.wikipedia.org/wiki/Theodore_W._Richards
Th�ophile Gautier	http://en.wikipedia.org/wiki/Th%E9ophile_Gautier
Theresa LePore	http://en.wikipedia.org/wiki/Theresa_LePore
Theresa May	http://en.wikipedia.org/wiki/Theresa_May
Theresa Russell	http://en.wikipedia.org/wiki/Theresa_Russell
Theresa Villiers	http://en.wikipedia.org/wiki/Theresa_Villiers
Therese Coffey	http://en.wikipedia.org/wiki/Therese_Coffey
Thierry Henry	http://en.wikipedia.org/wiki/Thierry_Henry
Thom Filicia	http://en.wikipedia.org/wiki/Thom_Filicia
Thom Gunn	http://en.wikipedia.org/wiki/Thom_Gunn
Thom Mayne	http://en.wikipedia.org/wiki/Thom_Mayne
Thom Yorke	http://en.wikipedia.org/wiki/Thom_Yorke
Thomas � Kempis	http://en.wikipedia.org/wiki/Thomas_%E0_Kempis
Thomas A. Luken	http://en.wikipedia.org/wiki/Thomas_A._Luken
Thomas A. Riggs	http://en.wikipedia.org/wiki/Thomas_Christmas_Riggs,_Jr.
Thomas Addison	http://en.wikipedia.org/wiki/Thomas_Addison
Thomas Allen	http://en.wikipedia.org/wiki/Tom_Allen_(comedian)
Thomas Andrews Hendricks	http://en.wikipedia.org/wiki/Thomas_Andrews_Hendricks
Thomas Arundel	http://en.wikipedia.org/wiki/Thomas_Arundel
Thomas B. Allen	http://en.wikipedia.org/wiki/Thomas_B._Allen_(author)
Thomas Babington Macaulay	http://en.wikipedia.org/wiki/Thomas_Babington_Macaulay
Thomas Bailey Aldrich	http://en.wikipedia.org/wiki/Thomas_Bailey_Aldrich
Thomas Becket	http://en.wikipedia.org/wiki/Thomas_Becket
Thomas Berger	http://en.wikipedia.org/wiki/Thomas_Berger_(novelist)
Thomas Bewick	http://en.wikipedia.org/wiki/Thomas_Bewick
Thomas Bilney	http://en.wikipedia.org/wiki/Thomas_Bilney
Thomas Bodley	http://en.wikipedia.org/wiki/Thomas_Bodley
Thomas Bulfinch	http://en.wikipedia.org/wiki/Thomas_Bulfinch
Thomas Burnet	http://en.wikipedia.org/wiki/Thomas_Burnet
Thomas C. Schelling	http://en.wikipedia.org/wiki/Thomas_C._Schelling
Thomas Cahill	http://en.wikipedia.org/wiki/Thomas_Cahill
Thomas Carew	http://en.wikipedia.org/wiki/Thomas_Carew
Thomas Carlyle	http://en.wikipedia.org/wiki/Thomas_Carlyle
Thomas Carper	http://en.wikipedia.org/wiki/Thomas_Carper
Thomas Cartwright	http://en.wikipedia.org/wiki/Thomas_Cartwright_(Puritan)
Thomas Cavanagh	http://en.wikipedia.org/wiki/Thomas_Cavanagh
Thomas Cavendish	http://en.wikipedia.org/wiki/Thomas_Cavendish
Thomas Chalmers	http://en.wikipedia.org/wiki/Thomas_Chalmers
Thomas Chatterton	http://en.wikipedia.org/wiki/Thomas_Chatterton
Thomas Cochrane	http://en.wikipedia.org/wiki/Thomas_Cochrane,_10th_Earl_of_Dundonald
Thomas Cole	http://en.wikipedia.org/wiki/Thomas_Cole
Thomas Cranmer	http://en.wikipedia.org/wiki/Thomas_Cranmer
Thomas Cromwell	http://en.wikipedia.org/wiki/Thomas_Cromwell
Thomas Dangerfield	http://en.wikipedia.org/wiki/Thomas_Dangerfield
Thomas Daschle	http://en.wikipedia.org/wiki/Thomas_Daschle
Thomas Davidson	http://en.wikipedia.org/wiki/Thomas_Davidson_(palaeontologist)
Thomas de Keyser	http://en.wikipedia.org/wiki/Thomas_de_Keyser
Thomas De Quincey	http://en.wikipedia.org/wiki/Thomas_De_Quincey
Thomas Dekker	http://en.wikipedia.org/wiki/Thomas_Dekker_(writer)
Thomas Dempster	http://en.wikipedia.org/wiki/Thomas_Dempster
Thomas Docherty	http://en.wikipedia.org/wiki/Thomas_Docherty_(politician)
Thomas Dolby	http://en.wikipedia.org/wiki/Thomas_Dolby
Thomas E. Dewey	http://en.wikipedia.org/wiki/Thomas_E._Dewey
Thomas E. Petri	http://en.wikipedia.org/wiki/Thomas_E._Petri
Thomas Eagleton	http://en.wikipedia.org/wiki/Thomas_Eagleton
Thomas Edison	http://en.wikipedia.org/wiki/Thomas_Edison
Thomas Erastus	http://en.wikipedia.org/wiki/Thomas_Erastus
Thomas Ewing	http://en.wikipedia.org/wiki/Thomas_Ewing
Thomas F. Eagleton	http://en.wikipedia.org/wiki/Thomas_F._Eagleton
Thomas F. Hartnett	http://en.wikipedia.org/wiki/Thomas_F._Hartnett
Thomas Fran�ois Burgers	http://en.wikipedia.org/wiki/Thomas_Fran%E7ois_Burgers
Thomas Frank	http://en.wikipedia.org/wiki/Thomas_Frank
Thomas Friedman	http://en.wikipedia.org/wiki/Thomas_Friedman
Thomas Frognall Dibdin	http://en.wikipedia.org/wiki/Thomas_Frognall_Dibdin
Thomas Gage	http://en.wikipedia.org/wiki/Thomas_Gage
Thomas Gainsborough	http://en.wikipedia.org/wiki/Thomas_Gainsborough
Thomas Gaisford	http://en.wikipedia.org/wiki/Thomas_Gaisford
Thomas Gibson	http://en.wikipedia.org/wiki/Thomas_Gibson
Thomas Gold	http://en.wikipedia.org/wiki/Thomas_Gold
Thomas Gray	http://en.wikipedia.org/wiki/Thomas_Gray
Thomas H. Cruikshank	http://en.wikipedia.org/wiki/Thomas_H._Cruikshank
Thomas H. Kean	http://en.wikipedia.org/wiki/Thomas_H._Kean
Thomas H. Kean, Jr.	http://en.wikipedia.org/wiki/Thomas_H._Kean%2C_Jr.
Thomas Haden Church	http://en.wikipedia.org/wiki/Thomas_Haden_Church
Thomas Hardy	http://en.wikipedia.org/wiki/Thomas_Hardy
Thomas Harris	http://en.wikipedia.org/wiki/Thomas_Harris
Thomas Hart Benton	http://en.wikipedia.org/wiki/Thomas_Hart_Benton_(painter)
Thomas Hart Benton	http://en.wikipedia.org/wiki/Thomas_Hart_Benton_(senator)
Thomas Hearne	http://en.wikipedia.org/wiki/Thomas_Hearne
Thomas Hearns	http://en.wikipedia.org/wiki/Thomas_Hearns
Thomas Henry Huxley	http://en.wikipedia.org/wiki/Thomas_Henry_Huxley
Thomas Heywood	http://en.wikipedia.org/wiki/Thomas_Heywood
Thomas Hobbes	http://en.wikipedia.org/wiki/Thomas_Hobbes
Thomas Holcroft	http://en.wikipedia.org/wiki/Thomas_Holcroft
Thomas Hood	http://en.wikipedia.org/wiki/Thomas_Hood
Thomas Hooker	http://en.wikipedia.org/wiki/Thomas_Hooker
Thomas Hughes	http://en.wikipedia.org/wiki/Thomas_Hughes
Thomas Hutchinson	http://en.wikipedia.org/wiki/Thomas_Hutchinson_(governor)
Thomas Ian Griffith	http://en.wikipedia.org/wiki/Thomas_Ian_Griffith
Thomas Ian Nicholas	http://en.wikipedia.org/wiki/Thomas_Ian_Nicholas
Thomas J. "Jerry" Huckaby	http://en.wikipedia.org/wiki/Jerry_Huckaby
Thomas J. Bliley, Jr.	http://en.wikipedia.org/wiki/Thomas_J._Bliley%2C_Jr.
Thomas J. Downey	http://en.wikipedia.org/wiki/Thomas_J._Downey
Thomas J. Falk	http://en.wikipedia.org/wiki/Thomas_J._Falk
Thomas J. Manton	http://en.wikipedia.org/wiki/Thomas_J._Manton
Thomas J. Usher	http://en.wikipedia.org/wiki/Thomas_Usher
Thomas J. Watson	http://en.wikipedia.org/wiki/Thomas_J._Watson
Thomas Jane	http://en.wikipedia.org/wiki/Thomas_Jane
Thomas Jefferson	http://en.wikipedia.org/wiki/Thomas_Jefferson
Thomas Keller	http://en.wikipedia.org/wiki/Thomas_Keller
Thomas Keneally	http://en.wikipedia.org/wiki/Thomas_Keneally
Thomas Killigrew	http://en.wikipedia.org/wiki/Thomas_Killigrew
Thomas King Forcade	http://en.wikipedia.org/wiki/Thomas_King_Forcade
Thomas Kinkade	http://en.wikipedia.org/wiki/Thomas_Kinkade
Thomas Klestil	http://en.wikipedia.org/wiki/Thomas_Klestil
Thomas Kuhn	http://en.wikipedia.org/wiki/Thomas_Kuhn
Thomas Kyd	http://en.wikipedia.org/wiki/Thomas_Kyd
Thomas Lennon	http://en.wikipedia.org/wiki/Thomas_Lennon_(actor)
Thomas Linacre	http://en.wikipedia.org/wiki/Thomas_Linacre
Thomas Love Peacock	http://en.wikipedia.org/wiki/Thomas_Love_Peacock
Thomas M. Foglietta	http://en.wikipedia.org/wiki/Thomas_M._Foglietta
Thomas M. Ryan	http://en.wikipedia.org/wiki/Thomas_Ryan_(businessman)
Thomas M. Siebel	http://en.wikipedia.org/wiki/Thomas_Siebel
Thomas Malthus	http://en.wikipedia.org/wiki/Thomas_Malthus
Thomas Mann	http://en.wikipedia.org/wiki/Thomas_Mann
Thomas May	http://en.wikipedia.org/wiki/Thomas_May
Thomas McGuane	http://en.wikipedia.org/wiki/Thomas_McGuane
Thomas Menino	http://en.wikipedia.org/wiki/Thomas_Menino
Thomas Merton	http://en.wikipedia.org/wiki/Thomas_Merton
Thomas Middleton	http://en.wikipedia.org/wiki/Thomas_Middleton
Thomas Mitchell	http://en.wikipedia.org/wiki/Thomas_Mitchell_(actor)
Thomas Monaghan	http://en.wikipedia.org/wiki/Tom_Monaghan
Thomas Morley	http://en.wikipedia.org/wiki/Thomas_Morley
Thomas Morton	http://en.wikipedia.org/wiki/Thomas_Morton_(colonist)
Thomas M�nzer	http://en.wikipedia.org/wiki/Thomas_M%FCnzer
Thomas N. Kindness	http://en.wikipedia.org/wiki/Thomas_N._Kindness
Thomas Nagel	http://en.wikipedia.org/wiki/Thomas_Nagel
Thomas Nashe	http://en.wikipedia.org/wiki/Thomas_Nashe
Thomas Nast	http://en.wikipedia.org/wiki/Thomas_Nast
Thomas Nelson Page	http://en.wikipedia.org/wiki/Thomas_Nelson_Page
Thomas Newcomen	http://en.wikipedia.org/wiki/Thomas_Newcomen
Thomas Otway	http://en.wikipedia.org/wiki/Thomas_Otway
Thomas P. O'Neill, Jr.	http://en.wikipedia.org/wiki/Thomas_P._O%27Neill%2C_Jr.
Thomas P. Stafford	http://en.wikipedia.org/wiki/Thomas_P._Stafford
Thomas Paine	http://en.wikipedia.org/wiki/Thomas_Paine
Thomas Parnell	http://en.wikipedia.org/wiki/Thomas_Parnell
Thomas Parr	http://en.wikipedia.org/wiki/Old_Tom_Parr
Thomas Penfield Jackson	http://en.wikipedia.org/wiki/Thomas_Penfield_Jackson
Thomas Percy	http://en.wikipedia.org/wiki/Thomas_Percy
Thomas Petri	http://en.wikipedia.org/wiki/Thomas_Petri
Thomas Pickering	http://en.wikipedia.org/wiki/Thomas_R._Pickering
Thomas Pinckney	http://en.wikipedia.org/wiki/Thomas_Pinckney
Thomas Pynchon	http://en.wikipedia.org/wiki/Thomas_Pynchon
Thomas R. Carper	http://en.wikipedia.org/wiki/Thomas_R._Carper
Thomas R. Cech	http://en.wikipedia.org/wiki/Thomas_R._Cech
Thomas R. Marshall	http://en.wikipedia.org/wiki/Thomas_R._Marshall
Thomas Reynolds	http://en.wikipedia.org/wiki/Thomas_Reynolds
Thomas Rowlandson	http://en.wikipedia.org/wiki/Thomas_Rowlandson
Thomas S. Foley	http://en.wikipedia.org/wiki/Thomas_S._Foley
Thomas S. Gates	http://en.wikipedia.org/wiki/Thomas_S._Gates
Thomas S. Kleppe	http://en.wikipedia.org/wiki/Thomas_S._Kleppe
Thomas Shadwell	http://en.wikipedia.org/wiki/Thomas_Shadwell
Thomas Sheraton	http://en.wikipedia.org/wiki/Thomas_Sheraton
Thomas Southerne	http://en.wikipedia.org/wiki/Thomas_Southerne
Thomas Sowell	http://en.wikipedia.org/wiki/Thomas_Sowell
Thomas Stothard	http://en.wikipedia.org/wiki/Thomas_Stothard
Thomas Stucley	http://en.wikipedia.org/wiki/Thomas_Stucley
Thomas Sully	http://en.wikipedia.org/wiki/Thomas_Sully
Thomas Sumter	http://en.wikipedia.org/wiki/Thomas_Sumter
Thomas Sydenham	http://en.wikipedia.org/wiki/Thomas_Sydenham
Thomas T. Noguchi	http://en.wikipedia.org/wiki/Thomas_Noguchi
Thomas Tallis	http://en.wikipedia.org/wiki/Thomas_Tallis
Thomas Telford	http://en.wikipedia.org/wiki/Thomas_Telford
Thomas Urquhart	http://en.wikipedia.org/wiki/Thomas_Urquhart
Thomas Vaughan	http://en.wikipedia.org/wiki/Thomas_Vaughan_(philosopher)
Thomas Vilsack	http://en.wikipedia.org/wiki/Thomas_Vilsack
Thomas Walsingham	http://en.wikipedia.org/wiki/Thomas_Walsingham
Thomas Warton	http://en.wikipedia.org/wiki/Thomas_Warton
Thomas Watson	http://en.wikipedia.org/wiki/Thomas_Watson_(poet)
Thomas Wolfe	http://en.wikipedia.org/wiki/Thomas_Wolfe
Thomas Wolsey	http://en.wikipedia.org/wiki/Thomas_Wolsey
Thor Heyerdahl	http://en.wikipedia.org/wiki/Thor_Heyerdahl
Thora Birch	http://en.wikipedia.org/wiki/Thora_Birch
Thora Hird	http://en.wikipedia.org/wiki/Thora_Hird
Thornton Wilder	http://en.wikipedia.org/wiki/Thornton_Wilder
Thorstein Veblen	http://en.wikipedia.org/wiki/Thorstein_Veblen
Thurgood Marshall	http://en.wikipedia.org/wiki/Thurgood_Marshall
Thurl Ravenscroft	http://en.wikipedia.org/wiki/Thurl_Ravenscroft
Thurlow Weed	http://en.wikipedia.org/wiki/Thurlow_Weed
Thurston Moore	http://en.wikipedia.org/wiki/Thurston_Moore
Tia Carrere	http://en.wikipedia.org/wiki/Tia_Carrere
Tia Mowry	http://en.wikipedia.org/wiki/Tia_Mowry
Tichina Arnold	http://en.wikipedia.org/wiki/Tichina_Arnold
Tiffani Amber Thiessen	http://en.wikipedia.org/wiki/Tiffani_Amber_Thiessen
Tiger Woods	http://en.wikipedia.org/wiki/Tiger_Woods
Tigran Sargsyan	http://en.wikipedia.org/wiki/Tigran_Sargsyan
Tiki Barber	http://en.wikipedia.org/wiki/Tiki_Barber
Tilda Swinton	http://en.wikipedia.org/wiki/Tilda_Swinton
Till Lindemann	http://en.wikipedia.org/wiki/Till_Lindemann
Tillie Olsen	http://en.wikipedia.org/wiki/Tillie_Olsen
Tillman Thomas	http://en.wikipedia.org/wiki/Tillman_Thomas
Tim Allen	http://en.wikipedia.org/wiki/Tim_Allen
Tim Armstrong	http://en.wikipedia.org/wiki/Tim_Armstrong
Tim Babcock	http://en.wikipedia.org/wiki/Tim_Babcock
Tim Berners-Lee	http://en.wikipedia.org/wiki/Tim_Berners-Lee
Tim Bray	http://en.wikipedia.org/wiki/Tim_Bray
Tim Buckley	http://en.wikipedia.org/wiki/Tim_Buckley
Tim Burton	http://en.wikipedia.org/wiki/Tim_Burton
Tim Considine	http://en.wikipedia.org/wiki/Tim_Considine
Tim Conway	http://en.wikipedia.org/wiki/Tim_Conway
Tim Curry	http://en.wikipedia.org/wiki/Tim_Curry
Tim DeLaughter	http://en.wikipedia.org/wiki/Tim_DeLaughter
Tim Duncan	http://en.wikipedia.org/wiki/Tim_Duncan
Tim Farron	http://en.wikipedia.org/wiki/Tim_Farron
Tim Finn	http://en.wikipedia.org/wiki/Tim_Finn
Tim Gane	http://en.wikipedia.org/wiki/Tim_Gane
Tim Holden	http://en.wikipedia.org/wiki/Tim_Holden
Tim Holt	http://en.wikipedia.org/wiki/Tim_Holt
Tim Hudson	http://en.wikipedia.org/wiki/Tim_Hudson
Tim Johnson	http://en.wikipedia.org/wiki/Tim_Johnson_(U.S._Representative)
Tim Johnson	http://en.wikipedia.org/wiki/Tim_Johnson_(U.S._Senator)
Tim Kaine	http://en.wikipedia.org/wiki/Tim_Kaine
Tim Kaine	http://en.wikipedia.org/wiki/Tim_Kaine
Tim Kazurinsky	http://en.wikipedia.org/wiki/Tim_Kazurinsky
Tim LaHaye	http://en.wikipedia.org/wiki/Tim_LaHaye
Tim Loughton	http://en.wikipedia.org/wiki/Tim_Loughton
Tim Matheson	http://en.wikipedia.org/wiki/Tim_Matheson
Tim McGraw	http://en.wikipedia.org/wiki/Tim_McGraw
Tim McInnerny	http://en.wikipedia.org/wiki/Tim_McInnerny
Tim Meadows	http://en.wikipedia.org/wiki/Tim_Meadows
Tim Murphy	http://en.wikipedia.org/wiki/Tim_Murphy_(congressman)
Tim O'Brien	http://en.wikipedia.org/wiki/Tim_O'Brien_(author)
Tim O'Reilly	http://en.wikipedia.org/wiki/Tim_O%27Reilly
Tim Pawlenty	http://en.wikipedia.org/wiki/Tim_Pawlenty
Tim Pigott-Smith	http://en.wikipedia.org/wiki/Tim_Pigott-Smith
Tim Prusmack	http://en.wikipedia.org/wiki/Tim_Prusmack
Tim Reid	http://en.wikipedia.org/wiki/Tim_Reid
Tim Rice	http://en.wikipedia.org/wiki/Tim_Rice
Tim Robbins	http://en.wikipedia.org/wiki/Tim_Robbins
Tim Roth	http://en.wikipedia.org/wiki/Tim_Roth
Tim Russert	http://en.wikipedia.org/wiki/Tim_Russert
Tim Ryan	http://en.wikipedia.org/wiki/Tim_Ryan
Tim Valentine	http://en.wikipedia.org/wiki/Tim_Valentine
Tim Walz	http://en.wikipedia.org/wiki/Tim_Walz
Tim Yeo	http://en.wikipedia.org/wiki/Tim_Yeo
Timothy Bishop	http://en.wikipedia.org/wiki/Timothy_Bishop
Timothy Bottoms	http://en.wikipedia.org/wiki/Timothy_Bottoms
Timothy Busfield	http://en.wikipedia.org/wiki/Timothy_Busfield
Timothy Dalton	http://en.wikipedia.org/wiki/Timothy_Dalton
Timothy Daly	http://en.wikipedia.org/wiki/Timothy_Daly
Timothy Donnelly	http://en.wikipedia.org/wiki/Timothy_Donnelly
Timothy Dwight	http://en.wikipedia.org/wiki/Timothy_Dwight_IV
Timothy E. Wirth	http://en.wikipedia.org/wiki/Timothy_E._Wirth
Timothy Flanigan	http://en.wikipedia.org/wiki/Timothy_Flanigan
Timothy Geithner	http://en.wikipedia.org/wiki/Timothy_Geithner
Timothy Hutton	http://en.wikipedia.org/wiki/Timothy_Hutton
Timothy J. Penny	http://en.wikipedia.org/wiki/Timothy_J._Penny
Timothy J. Roemer	http://en.wikipedia.org/wiki/Timothy_J._Roemer
Timothy Koogle	http://en.wikipedia.org/wiki/Timothy_Koogle
Timothy Leary	http://en.wikipedia.org/wiki/Timothy_Leary
Timothy M. Donahue	http://en.wikipedia.org/wiki/Timothy_Donahue
Timothy McVeigh	http://en.wikipedia.org/wiki/Timothy_McVeigh
Timothy Olyphant	http://en.wikipedia.org/wiki/Timothy_Olyphant
Timothy Spall	http://en.wikipedia.org/wiki/Timothy_Spall
Timothy Treadwell	http://en.wikipedia.org/wiki/Timothy_Treadwell
Timothy West	http://en.wikipedia.org/wiki/Timothy_West
Tina Brown	http://en.wikipedia.org/wiki/Tina_Brown
Tina Charles	http://en.wikipedia.org/wiki/Tina_Charles_(singer)
Tina Fey	http://en.wikipedia.org/wiki/Tina_Fey
Tina Landon	http://en.wikipedia.org/wiki/Tina_Landon
Tina Louise	http://en.wikipedia.org/wiki/Tina_Louise
Tina Majorino	http://en.wikipedia.org/wiki/Tina_Majorino
Tina Turner	http://en.wikipedia.org/wiki/Tina_Turner
Tina Weymouth	http://en.wikipedia.org/wiki/Tina_Weymouth
Tina Yothers	http://en.wikipedia.org/wiki/Tina_Yothers
Tino Martinez	http://en.wikipedia.org/wiki/Tino_Martinez
Tiny Tim	http://en.wikipedia.org/wiki/Tiny_Tim_(musician)
Tionne "T-Boz" Watkins	http://en.wikipedia.org/wiki/Tionne_%22T-Boz%22_Watkins
Tip O'Neill	http://en.wikipedia.org/wiki/Tip_O%27Neill
Tipper Gore	http://en.wikipedia.org/wiki/Tipper_Gore
Tippi Hedren	http://en.wikipedia.org/wiki/Tippi_Hedren
Tish Ambrose	http://en.wikipedia.org/wiki/Tish_Ambrose
Tisha Campbell	http://en.wikipedia.org/wiki/Tisha_Campbell
Tito Jackson	http://en.wikipedia.org/wiki/Tito_Jackson
Tito Puente	http://en.wikipedia.org/wiki/Tito_Puente
Titus Oates	http://en.wikipedia.org/wiki/Titus_Oates
Titus Welliver	http://en.wikipedia.org/wiki/Titus_Welliver
Tobe Hooper	http://en.wikipedia.org/wiki/Tobe_Hooper
Tobe Hooper	http://en.wikipedia.org/wiki/Tobe_Hooper
Tobey Maguire	http://en.wikipedia.org/wiki/Tobey_Maguire
Tobias Asser	http://en.wikipedia.org/wiki/Tobias_Asser
Tobias Ellwood	http://en.wikipedia.org/wiki/Tobias_Ellwood
Tobias Smollett	http://en.wikipedia.org/wiki/Tobias_Smollett
Tobias Wolff	http://en.wikipedia.org/wiki/Tobias_Wolff
Toby Amies	http://en.wikipedia.org/wiki/Toby_Amies
Toby Huss	http://en.wikipedia.org/wiki/Toby_Huss
Toby Keith	http://en.wikipedia.org/wiki/Toby_Keith
Toby Perkins	http://en.wikipedia.org/wiki/Toby_Perkins
Toby Roth	http://en.wikipedia.org/wiki/Toby_Roth
Toby Young	http://en.wikipedia.org/wiki/Toby_Young
Tod Browning	http://en.wikipedia.org/wiki/Tod_Browning
Todd Akin	http://en.wikipedia.org/wiki/Todd_Akin
Todd Allen	http://en.wikipedia.org/wiki/Todd_Allen
Todd Barry	http://en.wikipedia.org/wiki/Todd_Barry
Todd Bridges	http://en.wikipedia.org/wiki/Todd_Bridges
Todd Gitlin	http://en.wikipedia.org/wiki/Todd_Gitlin
Todd Haynes	http://en.wikipedia.org/wiki/Todd_Haynes
Todd Holoubek	http://en.wikipedia.org/wiki/Todd_Holoubek
Todd McFarlane	http://en.wikipedia.org/wiki/Todd_McFarlane
Todd Platts	http://en.wikipedia.org/wiki/Todd_Platts
Todd Rundgren	http://en.wikipedia.org/wiki/Todd_Rundgren
Todd Solondz	http://en.wikipedia.org/wiki/Todd_Solondz
Todd Tiahrt	http://en.wikipedia.org/wiki/Todd_Tiahrt
Todor Zhivkov	http://en.wikipedia.org/wiki/Todor_Zhivkov
Togiola Tulafono	http://en.wikipedia.org/wiki/Togiola_Tulafono
Togiola Tulafono	http://en.wikipedia.org/wiki/Togiola_Tulafono
Togiola Tulafono	http://en.wikipedia.org/wiki/Togiola_Tulafono
Togo West	http://en.wikipedia.org/wiki/Togo_West
Tom Allen	http://en.wikipedia.org/wiki/Tom_Allen
Tom Allen	http://en.wikipedia.org/wiki/Tom_Allen
Tom Amandes	http://en.wikipedia.org/wiki/Tom_Amandes
Tom Anderson	http://en.wikipedia.org/wiki/Tom_Anderson_(MySpace)
Tom Araya	http://en.wikipedia.org/wiki/Tom_Araya
Tom Arnold	http://en.wikipedia.org/wiki/Tom_Arnold_(actor)
Tom Atkins	http://en.wikipedia.org/wiki/Tom_Atkins_(actor)
Tom Baker	http://en.wikipedia.org/wiki/Tom_Baker
Tom Barrett	http://en.wikipedia.org/wiki/Tom_Barrett_(politician)
Tom Berenger	http://en.wikipedia.org/wiki/Tom_Berenger
Tom Bergeron	http://en.wikipedia.org/wiki/Tom_Bergeron
Tom Bevill	http://en.wikipedia.org/wiki/Tom_Bevill
Tom Blenkinsop	http://en.wikipedia.org/wiki/Tom_Blenkinsop
Tom Bodett	http://en.wikipedia.org/wiki/Tom_Bodett
Tom Bosley	http://en.wikipedia.org/wiki/Tom_Bosley
Tom Bradley	http://en.wikipedia.org/wiki/Tom_Bradley_(politician)
Tom Brady	http://en.wikipedia.org/wiki/Tom_Brady
Tom Brake	http://en.wikipedia.org/wiki/Tom_Brake
Tom Brokaw	http://en.wikipedia.org/wiki/Tom_Brokaw
Tom Clancy	http://en.wikipedia.org/wiki/Tom_Clancy
Tom Clarke	http://en.wikipedia.org/wiki/Tom_Clarke_(politician)
Tom Coburn	http://en.wikipedia.org/wiki/Tom_Coburn
Tom Cole	http://en.wikipedia.org/wiki/Tom_Cole
Tom Coleman	http://en.wikipedia.org/wiki/Tom_Coleman
Tom Conti	http://en.wikipedia.org/wiki/Tom_Conti
Tom Conway	http://en.wikipedia.org/wiki/Tom_Conway
Tom Cora	http://en.wikipedia.org/wiki/Tom_Cora
Tom Courtenay	http://en.wikipedia.org/wiki/Tom_Courtenay
Tom Cruise	http://en.wikipedia.org/wiki/Tom_Cruise
Tom Daschle	http://en.wikipedia.org/wiki/Tom_Daschle
Tom Davis	http://en.wikipedia.org/wiki/Thomas_M._Davis
Tom DeLay	http://en.wikipedia.org/wiki/Tom_DeLay
Tom DeLay	http://en.wikipedia.org/wiki/Tom_DeLay
Tom DeLonge	http://en.wikipedia.org/wiki/Tom_DeLonge
Tom Dooley	http://en.wikipedia.org/wiki/Thomas_Anthony_Dooley_III
Tom Feeney	http://en.wikipedia.org/wiki/Tom_Feeney
Tom Felton	http://en.wikipedia.org/wiki/Tom_Felton
Tom Flores	http://en.wikipedia.org/wiki/Tom_Flores
Tom Fogerty	http://en.wikipedia.org/wiki/Tom_Fogerty
Tom Foley	http://en.wikipedia.org/wiki/Tom_Foley
Tom Ford	http://en.wikipedia.org/wiki/Tom_Ford
Tom Gjelten	http://en.wikipedia.org/wiki/Tom_Gjelten
Tom Golisano	http://en.wikipedia.org/wiki/Tom_Golisano
Tom Greatrex	http://en.wikipedia.org/wiki/Tom_Greatrex
Tom Green	http://en.wikipedia.org/wiki/Tom_Green
Tom Hanks	http://en.wikipedia.org/wiki/Tom_Hanks
Tom Harkin	http://en.wikipedia.org/wiki/Tom_Harkin
Tom Harkin	http://en.wikipedia.org/wiki/Tom_Harkin
Tom Harris	http://en.wikipedia.org/wiki/Tom_Harris_(politician)
Tom Hayden	http://en.wikipedia.org/wiki/Tom_Hayden
Tom Herman	http://en.wikipedia.org/wiki/Tom_Herman
Tom Hicks	http://en.wikipedia.org/wiki/Tom_Hicks
Tom Houghton	http://en.wikipedia.org/wiki/Tom_Houghton
Tom Hulce	http://en.wikipedia.org/wiki/Tom_Hulce
Tom Jarriel	http://en.wikipedia.org/wiki/Tom_Jarriel
Tom Jenkinson	http://en.wikipedia.org/wiki/Tom_Jenkinson
Tom Jones	http://en.wikipedia.org/wiki/Tom_Jones_(singer)
Tom Joyner	http://en.wikipedia.org/wiki/Tom_Joyner
Tom Kenny	http://en.wikipedia.org/wiki/Tom_Kenny
Tom Landry	http://en.wikipedia.org/wiki/Tom_Landry
Tom Lantos	http://en.wikipedia.org/wiki/Tom_Lantos
Tom Lantos	http://en.wikipedia.org/wiki/Tom_Lantos
Tom Latham	http://en.wikipedia.org/wiki/Tom_Latham
Tom Laughlin	http://en.wikipedia.org/wiki/Tom_Laughlin
Tom Lehrer	http://en.wikipedia.org/wiki/Tom_Lehrer
Tom Lenk	http://en.wikipedia.org/wiki/Tom_Lenk
Tom Lewis	http://en.wikipedia.org/wiki/Tom_Lewis_(politician)
Tom Leykis	http://en.wikipedia.org/wiki/Tom_Leykis
Tom Loeffler	http://en.wikipedia.org/wiki/Tom_Loeffler
Tom McCamus	http://en.wikipedia.org/wiki/Tom_McCamus
Tom McClintock	http://en.wikipedia.org/wiki/Tom_McClintock
Tom Metzger	http://en.wikipedia.org/wiki/Tom_Metzger
Tom Mix	http://en.wikipedia.org/wiki/Tom_Mix
Tom Morello	http://en.wikipedia.org/wiki/Tom_Morello
Tom Osborne	http://en.wikipedia.org/wiki/Tom_Osborne
Tom Paxton	http://en.wikipedia.org/wiki/Tom_Paxton
Tom Periello	http://en.wikipedia.org/wiki/Tom_Periello
Tom Peters	http://en.wikipedia.org/wiki/Tom_Peters
Tom Petty	http://en.wikipedia.org/wiki/Tom_Petty
Tom Poston	http://en.wikipedia.org/wiki/Tom_Poston
Tom Price	http://en.wikipedia.org/wiki/Tom_Price_(U.S._politician)
Tom Ridge	http://en.wikipedia.org/wiki/Tom_Ridge
Tom Ridge	http://en.wikipedia.org/wiki/Tom_Ridge
Tom Robbins	http://en.wikipedia.org/wiki/Tom_Robbins
Tom Rooney	http://en.wikipedia.org/wiki/Tom_Rooney_(politician)
Tom Rowlands	http://en.wikipedia.org/wiki/Tom_Rowlands
Tom Savini	http://en.wikipedia.org/wiki/Tom_Savini
Tom Scholz	http://en.wikipedia.org/wiki/Tom_Scholz
Tom Scott	http://en.wikipedia.org/wiki/Tom_Scott_(musician)
Tom Seaver	http://en.wikipedia.org/wiki/Tom_Seaver
Tom Selleck	http://en.wikipedia.org/wiki/Tom_Selleck
Tom Shales	http://en.wikipedia.org/wiki/Tom_Shales
Tom Silva	http://en.wikipedia.org/wiki/Tom_Silva
Tom Sizemore	http://en.wikipedia.org/wiki/Tom_Sizemore
Tom Skerritt	http://en.wikipedia.org/wiki/Tom_Skerritt
Tom Sneddon	http://en.wikipedia.org/wiki/Tom_Sneddon
Tom Snyder	http://en.wikipedia.org/wiki/Tom_Snyder
Tom Stemberg	http://en.wikipedia.org/wiki/Thomas_G._Stemberg
Tom Stoppard	http://en.wikipedia.org/wiki/Tom_Stoppard
Tom T. Hall	http://en.wikipedia.org/wiki/Tom_T._Hall
Tom Tancredo	http://en.wikipedia.org/wiki/Tom_Tancredo
Tom Tauke	http://en.wikipedia.org/wiki/Tom_Tauke
Tom Tryon	http://en.wikipedia.org/wiki/Tom_Tryon
Tom Udall	http://en.wikipedia.org/wiki/Tom_Udall
Tom Verlaine	http://en.wikipedia.org/wiki/Tom_Verlaine
Tom Vilsack	http://en.wikipedia.org/wiki/Tom_Vilsack
Tom Waits	http://en.wikipedia.org/wiki/Tom_Waits
Tom Watson	http://en.wikipedia.org/wiki/Tom_Watson_(golfer)
Tom Watson	http://en.wikipedia.org/wiki/Tom_Watson_(politician)
Tom Welling	http://en.wikipedia.org/wiki/Tom_Welling
Tom Wilkinson	http://en.wikipedia.org/wiki/Tom_Wilkinson
Tom Wolfe	http://en.wikipedia.org/wiki/Tom_Wolfe
Tom Wopat	http://en.wikipedia.org/wiki/Tom_Wopat
Tomas Alfredson	http://en.wikipedia.org/wiki/Tomas_Alfredson
Tomas Masaryk	http://en.wikipedia.org/wiki/Tomas_Masaryk
Tomaso Albinoni	http://en.wikipedia.org/wiki/Tomaso_Albinoni
Tom� Vera Cruz	http://en.wikipedia.org/wiki/Tom%E9_Vera_Cruz
Tommaso Campanella	http://en.wikipedia.org/wiki/Tommaso_Campanella
Tommaso Grossi	http://en.wikipedia.org/wiki/Tommaso_Grossi
Tommy Allen	http://en.wikipedia.org/wiki/Tommy_Allen_%28speedway_rider%29
Tommy Ambrose	http://en.wikipedia.org/wiki/Tommy_Ambrose
Tommy Bond	http://en.wikipedia.org/wiki/Tommy_Bond
Tommy Chong	http://en.wikipedia.org/wiki/Tommy_Chong
Tommy Davidson	http://en.wikipedia.org/wiki/Tommy_Davidson
Tommy Dorsey	http://en.wikipedia.org/wiki/Tommy_Dorsey
Tommy F. Robinson	http://en.wikipedia.org/wiki/Tommy_F._Robinson
Tommy Flanagan	http://en.wikipedia.org/wiki/Tommy_Flanagan_(actor)
Tommy Franks	http://en.wikipedia.org/wiki/Tommy_Franks
Tommy Hilfiger	http://en.wikipedia.org/wiki/Tommy_Hilfiger
Tommy Kirk	http://en.wikipedia.org/wiki/Tommy_Kirk
Tommy Lasorda	http://en.wikipedia.org/wiki/Tommy_Lasorda
Tommy Lee	http://en.wikipedia.org/wiki/Tommy_Lee
Tommy Lee Jones	http://en.wikipedia.org/wiki/Tommy_Lee_Jones
Tommy Mottola	http://en.wikipedia.org/wiki/Tommy_Mottola
Tommy Noonan	http://en.wikipedia.org/wiki/Tommy_Noonan
Tommy Ramone	http://en.wikipedia.org/wiki/Tommy_Ramone
Tommy Remengesau	http://en.wikipedia.org/wiki/Tommy_Remengesau
Tommy Rettig	http://en.wikipedia.org/wiki/Tommy_Rettig
Tommy Shaw	http://en.wikipedia.org/wiki/Tommy_Shaw
Tommy Smothers	http://en.wikipedia.org/wiki/Tommy_Smothers
Tommy Thompson	http://en.wikipedia.org/wiki/Tommy_Thompson
Tommy Tune	http://en.wikipedia.org/wiki/Tommy_Tune
Tone Loc	http://en.wikipedia.org/wiki/Tone_Loc
Toni Braxton	http://en.wikipedia.org/wiki/Toni_Braxton
Toni Cade Bambara	http://en.wikipedia.org/wiki/Toni_Cade_Bambara
Toni Collette	http://en.wikipedia.org/wiki/Toni_Collette
Toni Morrison	http://en.wikipedia.org/wiki/Toni_Morrison
Toni Onley	http://en.wikipedia.org/wiki/Toni_Onley
Tony Allen	http://en.wikipedia.org/wiki/Tony_Allen_%28basketball%29
Tony Baldry	http://en.wikipedia.org/wiki/Tony_Baldry
Tony Banks	http://en.wikipedia.org/wiki/Tony_Banks_(musician)
Tony Benn	http://en.wikipedia.org/wiki/Tony_Benn
Tony Bennett	http://en.wikipedia.org/wiki/Tony_Bennett
Tony Bill	http://en.wikipedia.org/wiki/Tony_Bill
Tony Blair	http://en.wikipedia.org/wiki/Tony_Blair
Tony Blair	http://en.wikipedia.org/wiki/Tony_Blair
Tony Blankley	http://en.wikipedia.org/wiki/Tony_Blankley
Tony Brown	http://en.wikipedia.org/wiki/Tony_Brown_(journalist)
Tony Coelho	http://en.wikipedia.org/wiki/Tony_Coelho
Tony Conrad	http://en.wikipedia.org/wiki/Tony_Conrad
Tony Cunningham	http://en.wikipedia.org/wiki/Tony_Cunningham
Tony Curtis	http://en.wikipedia.org/wiki/Tony_Curtis
Tony Danza	http://en.wikipedia.org/wiki/Tony_Danza
Tony Dorsett	http://en.wikipedia.org/wiki/Tony_Dorsett
Tony Dow	http://en.wikipedia.org/wiki/Tony_Dow
Tony Dungy	http://en.wikipedia.org/wiki/Tony_Dungy
Tony Franciosa	http://en.wikipedia.org/wiki/Tony_Franciosa
Tony Goldwyn	http://en.wikipedia.org/wiki/Tony_Goldwyn
Tony Gwynn	http://en.wikipedia.org/wiki/Tony_Gwynn
Tony Hancock	http://en.wikipedia.org/wiki/Tony_Hancock
Tony Hawk	http://en.wikipedia.org/wiki/Tony_Hawk
Tony Hayward	http://en.wikipedia.org/wiki/Tony_Hayward
Tony Hillerman	http://en.wikipedia.org/wiki/Tony_Hillerman
Tony Horwitz	http://en.wikipedia.org/wiki/Tony_Horwitz
Tony Iommi	http://en.wikipedia.org/wiki/Tony_Iommi
Tony James	http://en.wikipedia.org/wiki/Tony_James
Tony Kornheiser	http://en.wikipedia.org/wiki/Tony_Kornheiser
Tony Kushner	http://en.wikipedia.org/wiki/Tony_Kushner
Tony LaRussa	http://en.wikipedia.org/wiki/Tony_LaRussa
Tony Levin	http://en.wikipedia.org/wiki/Tony_Levin
Tony Lloyd	http://en.wikipedia.org/wiki/Tony_Lloyd
Tony Lo Bianco	http://en.wikipedia.org/wiki/Tony_Lo_Bianco
Tony Martin	http://en.wikipedia.org/wiki/Tony_Martin_(musician)
Tony Martinez	http://en.wikipedia.org/wiki/Tony_Martinez
Tony Millionaire	http://en.wikipedia.org/wiki/Tony_Millionaire
Tony Orlando	http://en.wikipedia.org/wiki/Tony_Orlando
Tony Oxley	http://en.wikipedia.org/wiki/Tony_Oxley
Tony P. Hall	http://en.wikipedia.org/wiki/Tony_P._Hall
Tony Parker	http://en.wikipedia.org/wiki/Tony_Parker
Tony Perkins	http://en.wikipedia.org/wiki/Tony_Perkins_(politician)
Tony Randall	http://en.wikipedia.org/wiki/Tony_Randall
Tony Richardson	http://en.wikipedia.org/wiki/Tony_Richardson
Tony Robbins	http://en.wikipedia.org/wiki/Tony_Robbins
Tony Scott	http://en.wikipedia.org/wiki/Tony_Scott
Tony Shalhoub	http://en.wikipedia.org/wiki/Tony_Shalhoub
Tony Sirico	http://en.wikipedia.org/wiki/Tony_Sirico
Tony Snow	http://en.wikipedia.org/wiki/Tony_Snow
Tony Stewart	http://en.wikipedia.org/wiki/Tony_Stewart
Tony Visconti	http://en.wikipedia.org/wiki/Tony_Visconti
Tony Yayo	http://en.wikipedia.org/wiki/Tony_Yayo
Tonya Harding	http://en.wikipedia.org/wiki/Tonya_Harding
Tonya Kay	http://en.wikipedia.org/wiki/Tonya_Kay
Too Short	http://en.wikipedia.org/wiki/Too_Short
Tookie Williams	http://en.wikipedia.org/wiki/Tookie_Williams
Toomas Hendrik Ilves	http://en.wikipedia.org/wiki/Toomas_Hendrik_Ilves
Toots Thielemans	http://en.wikipedia.org/wiki/Toots_Thielemans
Topher Grace	http://en.wikipedia.org/wiki/Topher_Grace
Tor Johnson	http://en.wikipedia.org/wiki/Tor_Johnson
Tori Amos	http://en.wikipedia.org/wiki/Tori_Amos
Tori Spelling	http://en.wikipedia.org/wiki/Tori_Spelling
Torquato Tasso	http://en.wikipedia.org/wiki/Torquato_Tasso
Torrie Wilson	http://en.wikipedia.org/wiki/Torrie_Wilson
Toru Iwatani	http://en.wikipedia.org/wiki/Toru_Iwatani
Toshir� Mifune	http://en.wikipedia.org/wiki/Toshir%F4_Mifune
Toumani Diabat�	http://en.wikipedia.org/wiki/Toumani_Diabat%E9
Toussaint L'Ouverture	http://en.wikipedia.org/wiki/Toussaint_L%27Ouverture
Tracee Ellis Ross	http://en.wikipedia.org/wiki/Tracee_Ellis_Ross
Tracey Crouch	http://en.wikipedia.org/wiki/Tracey_Crouch
Tracey Gold	http://en.wikipedia.org/wiki/Tracey_Gold
Tracey Ullman	http://en.wikipedia.org/wiki/Tracey_Ullman
Tracey Walter	http://en.wikipedia.org/wiki/Tracey_Walter
Traci Bingham	http://en.wikipedia.org/wiki/Traci_Bingham
Tracy Chapman	http://en.wikipedia.org/wiki/Tracy_Chapman
Tracy Chevalier	http://en.wikipedia.org/wiki/Tracy_Chevalier
Tracy Kidder	http://en.wikipedia.org/wiki/Tracy_Kidder
Tracy McGrady	http://en.wikipedia.org/wiki/Tracy_McGrady
Tracy Morgan	http://en.wikipedia.org/wiki/Tracy_Morgan
Tracy Nelson	http://en.wikipedia.org/wiki/Tracy_Nelson_(actress)
Tracy Pollan	http://en.wikipedia.org/wiki/Tracy_Pollan
Tracy Scoggins	http://en.wikipedia.org/wiki/Tracy_Scoggins
Traian Basescu	http://en.wikipedia.org/wiki/Traian_Basescu
Trajano Boccalini	http://en.wikipedia.org/wiki/Trajano_Boccalini
Tran Duc Luong	http://en.wikipedia.org/wiki/Tran_Duc_Luong
Travis Barker	http://en.wikipedia.org/wiki/Travis_Barker
Travis Childers	http://en.wikipedia.org/wiki/Travis_Childers
Travis Davis	http://en.wikipedia.org/wiki/Travis_Davis
Travis Fimmel	http://en.wikipedia.org/wiki/Travis_Fimmel
Travis Tritt	http://en.wikipedia.org/wiki/Travis_Tritt
Traylor Howard	http://en.wikipedia.org/wiki/Traylor_Howard
Tre Cool	http://en.wikipedia.org/wiki/Tre_Cool
Treat Williams	http://en.wikipedia.org/wiki/Treat_Williams
Trent Ford	http://en.wikipedia.org/wiki/Trent_Ford
Trent Franks	http://en.wikipedia.org/wiki/Trent_Franks
Trent Lott	http://en.wikipedia.org/wiki/Trent_Lott
Trent Lott	http://en.wikipedia.org/wiki/Trent_Lott
Trent Reznor	http://en.wikipedia.org/wiki/Trent_Reznor
Tress MacNeille	http://en.wikipedia.org/wiki/Tress_MacNeille
Trevor Allen	http://en.wikipedia.org/wiki/Trevor_Allen
Trevor Bolder	http://en.wikipedia.org/wiki/Trevor_Bolder
Trevor Brown	http://en.wikipedia.org/wiki/Trevor_Brown
Trevor Dunn	http://en.wikipedia.org/wiki/Trevor_Dunn
Trevor Horn	http://en.wikipedia.org/wiki/Trevor_Horn
Trevor Howard	http://en.wikipedia.org/wiki/Trevor_Howard
Trevor Huddleston	http://en.wikipedia.org/wiki/Trevor_Huddleston
Trevor Nunn	http://en.wikipedia.org/wiki/Trevor_Nunn
Trevor Rabin	http://en.wikipedia.org/wiki/Trevor_Rabin
Trey Anastasio	http://en.wikipedia.org/wiki/Trey_Anastasio
Trey Parker	http://en.wikipedia.org/wiki/Trey_Parker
Trey Songz	http://en.wikipedia.org/wiki/Trey_Songz
Trey Spruance	http://en.wikipedia.org/wiki/Trey_Spruance
Tricia Nixon	http://en.wikipedia.org/wiki/Tricia_Nixon
Trick Daddy	http://en.wikipedia.org/wiki/Trick_Daddy
Trina McGee	http://en.wikipedia.org/wiki/Trina_McGee
Trina Schart Hyman	http://en.wikipedia.org/wiki/Trina_Schart_Hyman
Trini Lopez	http://en.wikipedia.org/wiki/Trini_Lopez
Trip Hawkins	http://en.wikipedia.org/wiki/Trip_Hawkins
Triple H	http://en.wikipedia.org/wiki/Triple_H
Tris Speaker	http://en.wikipedia.org/wiki/Tris_Speaker
Trish Stratus	http://en.wikipedia.org/wiki/Trish_Stratus
Trisha Goddard	http://en.wikipedia.org/wiki/Trisha_Goddard
Trisha Yearwood	http://en.wikipedia.org/wiki/Trisha_Yearwood
Trishelle Cannatella	http://en.wikipedia.org/wiki/Trishelle_Cannatella
Trista Rehn	http://en.wikipedia.org/wiki/Trista_Rehn
Tristan A. Farnon	http://en.wikipedia.org/wiki/Tristan_A._Farnon
Tristan Tzara	http://en.wikipedia.org/wiki/Tristan_Tzara
Tristram Hunt	http://en.wikipedia.org/wiki/Tristram_Hunt
Trofim Lysenko	http://en.wikipedia.org/wiki/Trofim_Lysenko
Troy Aikman	http://en.wikipedia.org/wiki/Troy_Aikman
Troy Donahue	http://en.wikipedia.org/wiki/Troy_Donahue
Troy Garity	http://en.wikipedia.org/wiki/Troy_Garity
Troy Miller	http://en.wikipedia.org/wiki/Troy_Miller
Troy Vincent	http://en.wikipedia.org/wiki/Troy_Vincent
Truman Capote	http://en.wikipedia.org/wiki/Truman_Capote
Trygve Gulbranssen	http://en.wikipedia.org/wiki/Trygve_Gulbranssen
Trygve Lie	http://en.wikipedia.org/wiki/Trygve_Lie
Tsakhiagiyn Elbegdorj	http://en.wikipedia.org/wiki/Tsakhiagiyn_Elbegdorj
Tsar Alexander I	http://en.wikipedia.org/wiki/Tsar_Alexander_I
Tsar Alexander II	http://en.wikipedia.org/wiki/Tsar_Alexander_II
Tsar Alexis	http://en.wikipedia.org/wiki/Tsar_Alexis
Tsar Ivan III	http://en.wikipedia.org/wiki/Ivan_III_of_Russia
Tsar Ivan V	http://en.wikipedia.org/wiki/Ivan_V_of_Russia
Tsar Ivan VI	http://en.wikipedia.org/wiki/Ivan_VI_of_Russia
Tsar Michael	http://en.wikipedia.org/wiki/Michael_I_of_Russia
Tsar Nicholas I	http://en.wikipedia.org/wiki/Tsar_Nicholas_I
Tsar Nicholas II	http://en.wikipedia.org/wiki/Tsar_Nicholas_II
Tsar Paul I	http://en.wikipedia.org/wiki/Paul_I_of_Russia
Tsar Peter II	http://en.wikipedia.org/wiki/Peter_II_of_Russia
Tsar Peter III	http://en.wikipedia.org/wiki/Tsar_Peter_III
Tsar Vasily III	http://en.wikipedia.org/wiki/Vasili_III_of_Russia
Tsung-Dao Lee	http://en.wikipedia.org/wiki/Tsung-Dao_Lee
Tuanku Syed Sirajuddin ibni al-Marhum Syed Putra Jamalullail	http://en.wikipedia.org/wiki/Tuanku_Syed_Sirajuddin_ibni_al-Marhum_Syed_Putra_Jamalullail
Tucker Carlson	http://en.wikipedia.org/wiki/Tucker_Carlson
Tuesday Weld	http://en.wikipedia.org/wiki/Tuesday_Weld
Tufuga Efi	http://en.wikipedia.org/wiki/Tufuga_Efi
Tug McGraw	http://en.wikipedia.org/wiki/Tug_McGraw
Tuila'epa Sailele Malielegaoi	http://en.wikipedia.org/wiki/Tuila%27epa_Sailele_Malielegaoi
Tullio Levi-Civita	http://en.wikipedia.org/wiki/Tullio_Levi-Civita
Tunde Adebimpe	http://en.wikipedia.org/wiki/Tunde_Adebimpe
Tupac Shakur	http://en.wikipedia.org/wiki/Tupac_Shakur
Tura Satana	http://en.wikipedia.org/wiki/Tura_Satana
Turgut �zal	http://en.wikipedia.org/wiki/Turgut_%D6zal
Twiggy Ramirez	http://en.wikipedia.org/wiki/Twiggy_Ramirez
Twyla Tharp	http://en.wikipedia.org/wiki/Twyla_Tharp
Ty Cobb	http://en.wikipedia.org/wiki/Ty_Cobb
Ty Hardin	http://en.wikipedia.org/wiki/Ty_Hardin
Ty Herndon	http://en.wikipedia.org/wiki/Ty_Herndon
Ty Longley	http://en.wikipedia.org/wiki/Ty_Longley
Ty Pennington	http://en.wikipedia.org/wiki/Ty_Pennington
Tycho Brahe	http://en.wikipedia.org/wiki/Tycho_Brahe
Tyler Christopher	http://en.wikipedia.org/wiki/Tyler_Christopher_(actor)
Tyler Florence	http://en.wikipedia.org/wiki/Tyler_Florence
Tyler Hilton	http://en.wikipedia.org/wiki/Tyler_Hilton
Tyler Hoechlin	http://en.wikipedia.org/wiki/Tyler_Hoechlin
Tyler Perry	http://en.wikipedia.org/wiki/Tyler_Perry
Tyne Daly	http://en.wikipedia.org/wiki/Tyne_Daly
Typhoid Mary	http://en.wikipedia.org/wiki/Typhoid_Mary
Tyra Banks	http://en.wikipedia.org/wiki/Tyra_Banks
Tyrees Allen	http://en.wikipedia.org/wiki/Tyrees_Allen
Tyrone Power	http://en.wikipedia.org/wiki/Tyrone_Power
Tyson Beckford	http://en.wikipedia.org/wiki/Tyson_Beckford
U Aung San	http://en.wikipedia.org/wiki/U_Aung_San
U Thant	http://en.wikipedia.org/wiki/U_Thant
Ub Iwerks	http://en.wikipedia.org/wiki/Ub_Iwerks
Uday Hussein	http://en.wikipedia.org/wiki/Uday_Hussein
Udo Kier	http://en.wikipedia.org/wiki/Udo_Kier
Ugo Foscolo	http://en.wikipedia.org/wiki/Ugo_Foscolo
Ulisse Aldrovandi	http://en.wikipedia.org/wiki/Ulisse_Aldrovandi
Ulrich von Hutten	http://en.wikipedia.org/wiki/Ulrich_von_Hutten
Ulysses S. Grant	http://en.wikipedia.org/wiki/Ulysses_S._Grant
Uma Thurman	http://en.wikipedia.org/wiki/Uma_Thurman
Umberto Boccioni	http://en.wikipedia.org/wiki/Umberto_Boccioni
Umberto Eco	http://en.wikipedia.org/wiki/Umberto_Eco
Uncle Kracker	http://en.wikipedia.org/wiki/Uncle_Kracker
Upton Sinclair	http://en.wikipedia.org/wiki/Upton_Sinclair
Uri Geller	http://en.wikipedia.org/wiki/Uri_Geller
Ursula Andress	http://en.wikipedia.org/wiki/Ursula_Andress
Ursula K. Le Guin	http://en.wikipedia.org/wiki/Ursula_K._Le_Guin
Uta Hagen	http://en.wikipedia.org/wiki/Uta_Hagen
Utada Hikaru	http://en.wikipedia.org/wiki/Utada_Hikaru
Uwe Boll	http://en.wikipedia.org/wiki/Uwe_Boll
V. C. Andrews	http://en.wikipedia.org/wiki/V._C._Andrews
V. S. Naipaul	http://en.wikipedia.org/wiki/V._S._Naipaul
V. S. Pritchett	http://en.wikipedia.org/wiki/V._S._Pritchett
Vachel Lindsay	http://en.wikipedia.org/wiki/Vachel_Lindsay
Vaclav Havel	http://en.wikipedia.org/wiki/Vaclav_Havel
Vaclav Klaus	http://en.wikipedia.org/wiki/Vaclav_Klaus
V�clav Klaus	http://en.wikipedia.org/wiki/V%E1clav_Klaus
Vaginal Davis 	http://en.wikipedia.org/wiki/Vaginal_Davis_
Vaira Vike-Freiberga	http://en.wikipedia.org/wiki/Vaira_Vike-Freiberga
Val Fitch	http://en.wikipedia.org/wiki/Val_Fitch
Val Guest	http://en.wikipedia.org/wiki/Val_Guest
Val Kilmer	http://en.wikipedia.org/wiki/Val_Kilmer
Valdas Adamkus	http://en.wikipedia.org/wiki/Valdas_Adamkus
Valdis Dombrovskis	http://en.wikipedia.org/wiki/Valdis_Dombrovskis
Valdis Zatlers	http://en.wikipedia.org/wiki/Valdis_Zatlers
Valentina Cortese	http://en.wikipedia.org/wiki/Valentina_Cortese
Valentino Rossi	http://en.wikipedia.org/wiki/Valentino_Rossi
Valeria Mazza	http://en.wikipedia.org/wiki/Valeria_Mazza
Valerie Bertinelli	http://en.wikipedia.org/wiki/Valerie_Bertinelli
Valerie Cruz	http://en.wikipedia.org/wiki/Valerie_Cruz
Valerie Harper	http://en.wikipedia.org/wiki/Valerie_Harper
Valerie Perrine	http://en.wikipedia.org/wiki/Valerie_Perrine
Valerie Plame	http://en.wikipedia.org/wiki/Valerie_Plame
Valerie Simpson	http://en.wikipedia.org/wiki/Valerie_Simpson
Valerie Solanas	http://en.wikipedia.org/wiki/Valerie_Solanas
Valerie Vaz	http://en.wikipedia.org/wiki/Valerie_Vaz
Val�ry Giscard d'Estaing	http://en.wikipedia.org/wiki/Val%E9ry_Giscard_d%27Estaing
Van Cliburn	http://en.wikipedia.org/wiki/Van_Cliburn
Van Heflin	http://en.wikipedia.org/wiki/Van_Heflin
Van Johnson	http://en.wikipedia.org/wiki/Van_Johnson
Van McCoy	http://en.wikipedia.org/wiki/Van_McCoy
Van Morrison	http://en.wikipedia.org/wiki/Van_Morrison
Van Williams	http://en.wikipedia.org/wiki/Van_Williams
Van Wyck Brooks	http://en.wikipedia.org/wiki/Van_Wyck_Brooks
Vance Amory	http://en.wikipedia.org/wiki/Vance_Amory
Vance Bourjaily	http://en.wikipedia.org/wiki/Vance_Bourjaily
Vance D. Coffman	http://en.wikipedia.org/wiki/Vance_D._Coffman
Vance Packard	http://en.wikipedia.org/wiki/Vance_Packard
Vanessa Amorosi	http://en.wikipedia.org/wiki/Vanessa_Amorosi
Vanessa Angel	http://en.wikipedia.org/wiki/Vanessa_Angel
Vanessa Carlton	http://en.wikipedia.org/wiki/Vanessa_Carlton
Vanessa Hudgens	http://en.wikipedia.org/wiki/Vanessa_Hudgens
Vanessa Incontrada	http://en.wikipedia.org/wiki/Vanessa_Incontrada
Vanessa Marcil	http://en.wikipedia.org/wiki/Vanessa_Marcil
Vanessa Paradis	http://en.wikipedia.org/wiki/Vanessa_Paradis
Vanessa Redgrave	http://en.wikipedia.org/wiki/Vanessa_Redgrave
Vanessa Williams	http://en.wikipedia.org/wiki/Vanessa_L._Williams
Vanilla Ice	http://en.wikipedia.org/wiki/Vanilla_Ice
Vanna White	http://en.wikipedia.org/wiki/Vanna_White
Vannevar Bush	http://en.wikipedia.org/wiki/Vannevar_Bush
Varg Vikernes	http://en.wikipedia.org/wiki/Varg_Vikernes
Vasco da Gama	http://en.wikipedia.org/wiki/Vasco_da_Gama
Vasco Nu�ez de Balboa	http://en.wikipedia.org/wiki/Vasco_Nu%F1ez_de_Balboa
Vasco Rossi	http://en.wikipedia.org/wiki/Vasco_Rossi
Vasile Tarlev	http://en.wikipedia.org/wiki/Vasile_Tarlev
Vaso Abashidze	http://en.wikipedia.org/wiki/Vaso_Abashidze
Vast Aire	http://en.wikipedia.org/wiki/Vast_Aire
Vaughan Kester	http://en.wikipedia.org/wiki/Vaughan_Kester
Ved Mehta	http://en.wikipedia.org/wiki/Ved_Mehta
Veit Stoss	http://en.wikipedia.org/wiki/Veit_Stoss
Velton Ray Bunch	http://en.wikipedia.org/wiki/Velton_Ray_Bunch
Vendela Kirsebom	http://en.wikipedia.org/wiki/Vendela_Kirsebom
Venerable Bede	http://en.wikipedia.org/wiki/Venerable_Bede
Venus Williams	http://en.wikipedia.org/wiki/Venus_Williams
Vera Alentova	http://en.wikipedia.org/wiki/Vera_Alentova
Vera Brittain	http://en.wikipedia.org/wiki/Vera_Brittain
Vera Lynn	http://en.wikipedia.org/wiki/Vera_Lynn
Vera Miles	http://en.wikipedia.org/wiki/Vera_Miles
Vera Ralston	http://en.wikipedia.org/wiki/Vera_Ralston
Vera Wang	http://en.wikipedia.org/wiki/Vera_Wang
Vern Yip	http://en.wikipedia.org/wiki/Vern_Yip
Verna Felton	http://en.wikipedia.org/wiki/Verna_Felton
Verne Lundquist	http://en.wikipedia.org/wiki/Verne_Lundquist
Verne Meisner	http://en.wikipedia.org/wiki/Verne_Meisner
Verne Troyer	http://en.wikipedia.org/wiki/Verne_Troyer
Vernon Bartlett	http://en.wikipedia.org/wiki/Vernon_Bartlett
Vernon Coaker	http://en.wikipedia.org/wiki/Vernon_Coaker
Vernon Ehlers	http://en.wikipedia.org/wiki/Vernon_Ehlers
Vernon Jordan	http://en.wikipedia.org/wiki/Vernon_Jordan
Vernon Louis Parrington	http://en.wikipedia.org/wiki/Vernon_Louis_Parrington
Vernon Sewell	http://en.wikipedia.org/wiki/Vernon_Sewell
Vernon Walters	http://en.wikipedia.org/wiki/Vernon_Walters
Vernor Vinge	http://en.wikipedia.org/wiki/Vernor_Vinge
Verona Feldbusch	http://en.wikipedia.org/wiki/Verona_Feldbusch
Veronica Cartwright	http://en.wikipedia.org/wiki/Veronica_Cartwright
Veronica Hamel	http://en.wikipedia.org/wiki/Veronica_Hamel
Veronica Lake	http://en.wikipedia.org/wiki/Veronica_Lake
Veronica Webb	http://en.wikipedia.org/wiki/Veronica_Webb
Vic Damone	http://en.wikipedia.org/wiki/Vic_Damone
Vic Dana	http://en.wikipedia.org/wiki/Vic_Dana
Vic Fazio	http://en.wikipedia.org/wiki/Vic_Fazio
Vic Morrow	http://en.wikipedia.org/wiki/Vic_Morrow
Vic Snyder	http://en.wikipedia.org/wiki/Vic_Snyder
Vic Tayback	http://en.wikipedia.org/wiki/Vic_Tayback
Vicente Fernandez	http://en.wikipedia.org/wiki/Vicente_Fernandez
Vicente Fox	http://en.wikipedia.org/wiki/Vicente_Fox
Vicente Fox	http://en.wikipedia.org/wiki/Vicente_Fox
Vicki Baum	http://en.wikipedia.org/wiki/Vicki_Baum
Vicki Lawrence	http://en.wikipedia.org/wiki/Vicki_Lawrence
Vicki Lewis	http://en.wikipedia.org/wiki/Vicki_Lewis
Vicki Mabrey	http://en.wikipedia.org/wiki/Vicki_Mabrey
Vicki Peterson	http://en.wikipedia.org/wiki/Vicki_Peterson
Vicky Botwright	http://en.wikipedia.org/wiki/Vicky_Botwright
Victor Argo	http://en.wikipedia.org/wiki/Victor_Argo
Victor Borge	http://en.wikipedia.org/wiki/Victor_Borge
Victor Buono	http://en.wikipedia.org/wiki/Victor_Buono
Victor Davis Hanson	http://en.wikipedia.org/wiki/Victor_Davis_Hanson
Victor de Laprade	http://en.wikipedia.org/wiki/Victor_de_Laprade
Victor Emmanuel II	http://en.wikipedia.org/wiki/Victor_Emmanuel_II
Victor Fleming	http://en.wikipedia.org/wiki/Victor_Fleming
Victor Francen	http://en.wikipedia.org/wiki/Victor_Francen
Victor Francis Hess	http://en.wikipedia.org/wiki/Victor_Francis_Hess
Victor French	http://en.wikipedia.org/wiki/Victor_French
Victor Garber	http://en.wikipedia.org/wiki/Victor_Garber
Victor Grignard	http://en.wikipedia.org/wiki/Victor_Grignard
Victor Horta	http://en.wikipedia.org/wiki/Victor_Horta
Victor Hugo	http://en.wikipedia.org/wiki/Victor_Hugo
Victor Jory	http://en.wikipedia.org/wiki/Victor_Jory
Victor Kiam	http://en.wikipedia.org/wiki/Victor_Kiam
Victor Krummenacher	http://en.wikipedia.org/wiki/Victor_Krummenacher
Victor Mature	http://en.wikipedia.org/wiki/Victor_Mature
Victor McLaglen	http://en.wikipedia.org/wiki/Victor_McLaglen
Victor Salva	http://en.wikipedia.org/wiki/Victor_Salva
Victor Sen Yung	http://en.wikipedia.org/wiki/Victor_Sen_Yung
Victor W. Turner	http://en.wikipedia.org/wiki/Victor_W._Turner
Victor Weisskopf	http://en.wikipedia.org/wiki/Victor_Weisskopf
Victor Willis	http://en.wikipedia.org/wiki/Victor_Willis
Victor Wong	http://en.wikipedia.org/wiki/Victor_Wong
Victor Young	http://en.wikipedia.org/wiki/Victor_Young
Victor Yushchenko	http://en.wikipedia.org/wiki/Victor_Yushchenko
Victoria Adams	http://en.wikipedia.org/wiki/Victoria_Beckham
Victoria Gotti	http://en.wikipedia.org/wiki/Victoria_Gotti
Victoria Jackson	http://en.wikipedia.org/wiki/Victoria_Jackson
Victoria Principal	http://en.wikipedia.org/wiki/Victoria_Principal
Victoria Rowell	http://en.wikipedia.org/wiki/Victoria_Rowell
Victoria Silvstedt	http://en.wikipedia.org/wiki/Victoria_Silvstedt
Victoria Toensing	http://en.wikipedia.org/wiki/Victoria_Toensing
Victorien Sardou	http://en.wikipedia.org/wiki/Victorien_Sardou
Vida Blue	http://en.wikipedia.org/wiki/Vida_Blue
Vida Guerra	http://en.wikipedia.org/wiki/Vida_Guerra
Vidal Sassoon	http://en.wikipedia.org/wiki/Vidal_Sassoon
Vidkun Quisling	http://en.wikipedia.org/wiki/Vidkun_Quisling
Viet Dinh	http://en.wikipedia.org/wiki/Viet_Dinh
Viggo Mortensen	http://en.wikipedia.org/wiki/Viggo_Mortensen
Vijay Singh	http://en.wikipedia.org/wiki/Vijay_Singh
Vikki Carr	http://en.wikipedia.org/wiki/Vikki_Carr
Viktor Chernomyrdin	http://en.wikipedia.org/wiki/Viktor_Chernomyrdin
Viktor Orb�n	http://en.wikipedia.org/wiki/Viktor_Orb%E1n
Viktor Yanukovych	http://en.wikipedia.org/wiki/Viktor_Yanukovych
Viktor Yushchenko	http://en.wikipedia.org/wiki/Viktor_Yushchenko
Ville Valo	http://en.wikipedia.org/wiki/Ville_Valo
Vin Diesel	http://en.wikipedia.org/wiki/Vin_Diesel
Vin Scully	http://en.wikipedia.org/wiki/Vin_Scully
Vin Weber	http://en.wikipedia.org/wiki/Vin_Weber
Vince Cable	http://en.wikipedia.org/wiki/Vince_Cable
Vince Carter	http://en.wikipedia.org/wiki/Vince_Carter
Vince Clarke	http://en.wikipedia.org/wiki/Vince_Clarke
Vince Edwards	http://en.wikipedia.org/wiki/Vince_Edwards
Vince Flynn	http://en.wikipedia.org/wiki/Vince_Flynn
Vince Foster	http://en.wikipedia.org/wiki/Vince_Foster
Vince Gill	http://en.wikipedia.org/wiki/Vince_Gill
Vince Lombardi	http://en.wikipedia.org/wiki/Vince_Lombardi
Vince McMahon	http://en.wikipedia.org/wiki/Vince_McMahon
Vince McMahon, Sr.	http://en.wikipedia.org/wiki/Vince_McMahon%2C_Sr.
Vince Neil	http://en.wikipedia.org/wiki/Vince_Neil
Vince Vaughn	http://en.wikipedia.org/wiki/Vince_Vaughn
Vincent Bugliosi	http://en.wikipedia.org/wiki/Vincent_Bugliosi
Vincent Cassel	http://en.wikipedia.org/wiki/Vincent_Cassel
Vincent Crane	http://en.wikipedia.org/wiki/Vincent_Crane
Vincent d'Indy	http://en.wikipedia.org/wiki/Vincent_d%27Indy
Vincent D'Onofrio	http://en.wikipedia.org/wiki/Vincent_D%27Onofrio
Vincent du Vigneaud	http://en.wikipedia.org/wiki/Vincent_du_Vigneaud
Vincent Gallo	http://en.wikipedia.org/wiki/Vincent_Gallo
Vincent Gardenia	http://en.wikipedia.org/wiki/Vincent_Gardenia
Vincent Gigante	http://en.wikipedia.org/wiki/Vincent_Gigante
Vincent Kartheiser	http://en.wikipedia.org/wiki/Vincent_Kartheiser
Vincent Margera	http://en.wikipedia.org/wiki/Vincent_Margera
Vincent Pastore	http://en.wikipedia.org/wiki/Vincent_Pastore
Vincent Perez	http://en.wikipedia.org/wiki/Vincent_Perez
Vincent Price	http://en.wikipedia.org/wiki/Vincent_Price
Vincent Schiavelli	http://en.wikipedia.org/wiki/Vincent_Schiavelli
Vincent Sherman	http://en.wikipedia.org/wiki/Vincent_Sherman
Vincent Spano	http://en.wikipedia.org/wiki/Vincent_Spano
Vincent van Gogh	http://en.wikipedia.org/wiki/Vincent_van_Gogh
Vincente Minnelli	http://en.wikipedia.org/wiki/Vincente_Minnelli
Vincenzo Bellini	http://en.wikipedia.org/wiki/Vincenzo_Bellini
Vincenzo Gioberti	http://en.wikipedia.org/wiki/Vincenzo_Gioberti
Ving Rhames	http://en.wikipedia.org/wiki/Ving_Rhames
Vinko Bogataj	http://en.wikipedia.org/wiki/Vinko_Bogataj
Vinnie Jones	http://en.wikipedia.org/wiki/Vinnie_Jones
Vinnie Paul	http://en.wikipedia.org/wiki/Vinnie_Paul
Vinnie Vincent	http://en.wikipedia.org/wiki/Vinnie_Vincent
Vinny Appice	http://en.wikipedia.org/wiki/Vinny_Appice
Vinny Testaverde	http://en.wikipedia.org/wiki/Vinny_Testaverde
Vint Cerf	http://en.wikipedia.org/wiki/Vint_Cerf
Viola Allen	http://en.wikipedia.org/wiki/Viola_Allen
Violent J	http://en.wikipedia.org/wiki/Violent_J
Violetta Chamorro	http://en.wikipedia.org/wiki/Violetta_Chamorro
Virender Sehwag	http://en.wikipedia.org/wiki/Virender_Sehwag
Virendra Sharma	http://en.wikipedia.org/wiki/Virendra_Sharma
Virgil Goode	http://en.wikipedia.org/wiki/Virgil_Goode
Virgil Thomson	http://en.wikipedia.org/wiki/Virgil_Thomson
Virgin Mary	http://en.wikipedia.org/wiki/Virgin_Mary
Virginia Christine	http://en.wikipedia.org/wiki/Virginia_Christine
Virginia Foxx	http://en.wikipedia.org/wiki/Virginia_Foxx
Virginia Madsen	http://en.wikipedia.org/wiki/Virginia_Madsen
Virginia Mayo	http://en.wikipedia.org/wiki/Virginia_Mayo
Virginia Smith	http://en.wikipedia.org/wiki/Virginia_Smith
Virginia Woolf	http://en.wikipedia.org/wiki/Virginia_Woolf
Virginie Ledoyen	http://en.wikipedia.org/wiki/Virginie_Ledoyen
Vitaly L. Ginzburg	http://en.wikipedia.org/wiki/Vitaly_L._Ginzburg
Vitas Gerulaitis	http://en.wikipedia.org/wiki/Vitas_Gerulaitis
Vito Fossella	http://en.wikipedia.org/wiki/Vito_Fossella
Vito Genovese	http://en.wikipedia.org/wiki/Vito_Genovese
Vittorio De Sica	http://en.wikipedia.org/wiki/Vittorio_De_Sica
Vitus Bering	http://en.wikipedia.org/wiki/Vitus_Bering
Viveca Novak	http://en.wikipedia.org/wiki/Viveca_Novak
Vivian Campbell	http://en.wikipedia.org/wiki/Vivian_Campbell
Vivian Richards	http://en.wikipedia.org/wiki/Vivian_Richards
Vivian Stanshall	http://en.wikipedia.org/wiki/Vivian_Stanshall
Vivian Vance	http://en.wikipedia.org/wiki/Vivian_Vance
Vivica Fox	http://en.wikipedia.org/wiki/Vivica_Fox
Vivien Leigh	http://en.wikipedia.org/wiki/Vivien_Leigh
Vivienne Westwood	http://en.wikipedia.org/wiki/Vivienne_Westwood
Vlad Filat	http://en.wikipedia.org/wiki/Vlad_Filat
Vlad the Impaler	http://en.wikipedia.org/wiki/Vlad_the_Impaler
Vladimir Arutyunian	http://en.wikipedia.org/wiki/Vladimir_Arutyunian
Vladimir Horowitz	http://en.wikipedia.org/wiki/Vladimir_Horowitz
Vladimir Komarov	http://en.wikipedia.org/wiki/Vladimir_Komarov
Vladimir Kramnik	http://en.wikipedia.org/wiki/Vladimir_Kramnik
Vladimir Nabokov	http://en.wikipedia.org/wiki/Vladimir_Nabokov
Vladimir Peniakoff	http://en.wikipedia.org/wiki/Vladimir_Peniakoff
Vladimir Prelog	http://en.wikipedia.org/wiki/Vladimir_Prelog
Vladimir Putin	http://en.wikipedia.org/wiki/Vladimir_Putin
Vladimir Sorokin	http://en.wikipedia.org/wiki/Vladimir_Sorokin
Vladimir Tatlin	http://en.wikipedia.org/wiki/Vladimir_Tatlin
Vladimir Voronin	http://en.wikipedia.org/wiki/Vladimir_Voronin
Vladimir Zhirinovsky	http://en.wikipedia.org/wiki/Vladimir_Zhirinovsky
Vlado Buckovski	http://en.wikipedia.org/wiki/Vlado_Buckovski
Vojislav Ko�tunica	http://en.wikipedia.org/wiki/Vojislav_Ko%9Atunica
Vojislav Seselj	http://en.wikipedia.org/wiki/Vojislav_Seselj
Volker Kriegel	http://en.wikipedia.org/wiki/Volker_Kriegel
Vsevolod Pudovkin	http://en.wikipedia.org/wiki/Vsevolod_Pudovkin
Vyacheslav Molotov	http://en.wikipedia.org/wiki/Vyacheslav_Molotov
W. Averell Harriman	http://en.wikipedia.org/wiki/W._Averell_Harriman
W. B. Maxwell	http://en.wikipedia.org/wiki/W._B._Maxwell
W. C. Fields	http://en.wikipedia.org/wiki/W._C._Fields
W. C. Handy	http://en.wikipedia.org/wiki/W._C._Handy
W. C. Wentworth	http://en.wikipedia.org/wiki/W._C._Wentworth
W. D. Snodgrass	http://en.wikipedia.org/wiki/W._D._Snodgrass
W. E. B. Du Bois	http://en.wikipedia.org/wiki/W._E._B._Du_Bois
W. Earl Brown	http://en.wikipedia.org/wiki/W._Earl_Brown
W. H. Auden	http://en.wikipedia.org/wiki/W._H._Auden
W. H. Hudson	http://en.wikipedia.org/wiki/W._H._Hudson
W. Henson Moore III	http://en.wikipedia.org/wiki/W._Henson_Moore_III
W. J. Usery	http://en.wikipedia.org/wiki/W._J._Usery
W. James McNerney Jr.	http://en.wikipedia.org/wiki/W._James_McNerney_Jr.
W. Mark Felt	http://en.wikipedia.org/wiki/W._Mark_Felt
W. Michael Blumenthal	http://en.wikipedia.org/wiki/W._Michael_Blumenthal
W. Richard Stevens	http://en.wikipedia.org/wiki/W._Richard_Stevens
W. S. Gilbert	http://en.wikipedia.org/wiki/W._S._Gilbert
W. S. Merwin	http://en.wikipedia.org/wiki/W._S._Merwin
W. S. Van Dyke	http://en.wikipedia.org/wiki/W._S._Van_Dyke
W. Somerset Maugham	http://en.wikipedia.org/wiki/W._Somerset_Maugham
W. W. Jacobs	http://en.wikipedia.org/wiki/W._W._Jacobs
W.D. Amaradeva	http://en.wikipedia.org/wiki/W.D._Amaradeva
W.V. Grant, Jr.	http://en.wikipedia.org/wiki/W._V._Grant
Waclaw Sierpinski	http://en.wikipedia.org/wiki/Waclaw_Sierpinski
Wade Boggs	http://en.wikipedia.org/wiki/Wade_Boggs
Wade Hampton	http://en.wikipedia.org/wiki/Wade_Hampton_III
Walafrid Strabo	http://en.wikipedia.org/wiki/Walafrid_Strabo
Walid Jumblatt	http://en.wikipedia.org/wiki/Walid_Jumblatt
Walker Percy	http://en.wikipedia.org/wiki/Walker_Percy
Wallace Beery	http://en.wikipedia.org/wiki/Wallace_Beery
Wallace Ford	http://en.wikipedia.org/wiki/Wallace_Ford
Wallace H. White, Jr.	http://en.wikipedia.org/wiki/Wallace_H._White%2C_Jr.
Wallace Hume Carothers	http://en.wikipedia.org/wiki/Wallace_Hume_Carothers
Wallace Langham	http://en.wikipedia.org/wiki/Wallace_Langham
Wallace Reid	http://en.wikipedia.org/wiki/Wallace_Reid
Wallace Shawn	http://en.wikipedia.org/wiki/Wallace_Shawn
Wallace Stegner	http://en.wikipedia.org/wiki/Wallace_Stegner
Wallace Stevens	http://en.wikipedia.org/wiki/Wallace_Stevens
Wallace Thurman	http://en.wikipedia.org/wiki/Wallace_Thurman
Wallis Simpson	http://en.wikipedia.org/wiki/Wallis_Simpson
Wally Cox	http://en.wikipedia.org/wiki/Wally_Cox
Wally George	http://en.wikipedia.org/wiki/Wally_George
Wally Herger	http://en.wikipedia.org/wiki/Wally_Herger
Wally O'Dell	http://en.wikipedia.org/wiki/Wally_O%27Dell
Wally Schirra	http://en.wikipedia.org/wiki/Wally_Schirra
Walt Disney	http://en.wikipedia.org/wiki/Walt_Disney
Walt Frazier	http://en.wikipedia.org/wiki/Walt_Frazier
Walt Hazzard	http://en.wikipedia.org/wiki/Walt_Hazzard
Walt Kelly	http://en.wikipedia.org/wiki/Walt_Kelly
Walt Rostow	http://en.wikipedia.org/wiki/Walt_Rostow
Walt Whitman	http://en.wikipedia.org/wiki/Walt_Whitman
Walter Abish	http://en.wikipedia.org/wiki/Walter_Abish
Walter Allen	http://en.wikipedia.org/wiki/Walter_Allen
Walter Annenberg	http://en.wikipedia.org/wiki/Walter_Annenberg
Walter B. Jones	http://en.wikipedia.org/wiki/Walter_B._Jones
Walter Baade	http://en.wikipedia.org/wiki/Walter_Baade
Walter Bagehot	http://en.wikipedia.org/wiki/Walter_Bagehot
Walter Beaman Jones, Sr.	http://en.wikipedia.org/wiki/Walter_Beaman_Jones%2C_Sr.
Walter Becker	http://en.wikipedia.org/wiki/Walter_Becker
Walter Bedell Smith	http://en.wikipedia.org/wiki/Walter_Bedell_Smith
Walter Benjamin	http://en.wikipedia.org/wiki/Walter_Benjamin
Walter Boughton Pitkin	http://en.wikipedia.org/wiki/Walter_Boughton_Pitkin
Walter Brennan	http://en.wikipedia.org/wiki/Walter_Brennan
Walter Crane	http://en.wikipedia.org/wiki/Walter_Crane
Walter Cronkite	http://en.wikipedia.org/wiki/Walter_Cronkite
Walter de la Mare	http://en.wikipedia.org/wiki/Walter_de_la_Mare
Walter Dean Burnham	http://en.wikipedia.org/wiki/Walter_Dean_Burnham
Walter E. Clark	http://en.wikipedia.org/wiki/Walter_Eli_Clark
Walter E. Fauntroy	http://en.wikipedia.org/wiki/Walter_E._Fauntroy
Walter E. Massey	http://en.wikipedia.org/wiki/Walter_E._Massey
Walter Gilbert	http://en.wikipedia.org/wiki/Walter_Gilbert
Walter Gropius	http://en.wikipedia.org/wiki/Walter_Gropius
Walter H. Brattain	http://en.wikipedia.org/wiki/Walter_H._Brattain
Walter Hagen	http://en.wikipedia.org/wiki/Walter_Hagen
Walter Hill	http://en.wikipedia.org/wiki/Walter_Hill_(filmmaker)
Walter Huston	http://en.wikipedia.org/wiki/Walter_Huston
Walter Isaacson	http://en.wikipedia.org/wiki/Walter_Isaacson
Walter J. Hickel	http://en.wikipedia.org/wiki/Walter_J._Hickel
Walter Johnson	http://en.wikipedia.org/wiki/Walter_Johnson
Walter Jon Williams	http://en.wikipedia.org/wiki/Walter_Jon_Williams
Walter Kerr	http://en.wikipedia.org/wiki/Walter_Kerr
Walter Knott	http://en.wikipedia.org/wiki/Walter_Knott
Walter Koenig	http://en.wikipedia.org/wiki/Walter_Koenig
Walter Kohn	http://en.wikipedia.org/wiki/Walter_Kohn
Walter Lang	http://en.wikipedia.org/wiki/Walter_Lang
Walter Leaf	http://en.wikipedia.org/wiki/Walter_Leaf
Walter Lippmann	http://en.wikipedia.org/wiki/Walter_Lippmann
Walter M. Miller, Jr.	http://en.wikipedia.org/wiki/Walter_M._Miller%2C_Jr.
Walter Macken	http://en.wikipedia.org/wiki/Walter_Macken
Walter Matthau	http://en.wikipedia.org/wiki/Walter_Matthau
Walter Mercado	http://en.wikipedia.org/wiki/Walter_Mercado
Walter Minnick	http://en.wikipedia.org/wiki/Walter_Minnick
Walter Mondale	http://en.wikipedia.org/wiki/Walter_Mondale
Walter Mosley	http://en.wikipedia.org/wiki/Walter_Mosley
Walter Mossberg	http://en.wikipedia.org/wiki/Walter_Mossberg
Walter P. Chrysler	http://en.wikipedia.org/wiki/Walter_P._Chrysler
Walter Pater	http://en.wikipedia.org/wiki/Walter_Pater
Walter Payton	http://en.wikipedia.org/wiki/Walter_Payton
Walter Pidgeon	http://en.wikipedia.org/wiki/Walter_Pidgeon
Walter Pincus	http://en.wikipedia.org/wiki/Walter_Pincus
Walter Piston	http://en.wikipedia.org/wiki/Walter_Piston
Walter Q. Gresham	http://en.wikipedia.org/wiki/Walter_Q._Gresham
Walter Reed	http://en.wikipedia.org/wiki/Walter_Reed
Walter Reuther	http://en.wikipedia.org/wiki/Walter_Reuther
Walter Russell Mead	http://en.wikipedia.org/wiki/Walter_Russell_Mead
Walter S. Carpenter, Jr.	http://en.wikipedia.org/wiki/Walter_S._Carpenter%2C_Jr.
Walter Salles	http://en.wikipedia.org/wiki/Walter_Salles
Walter Scheel	http://en.wikipedia.org/wiki/Walter_Scheel
Walter Slezak	http://en.wikipedia.org/wiki/Walter_Slezak
Walter Stoessel	http://en.wikipedia.org/wiki/Walter_Stoessel
Walter Ulbricht	http://en.wikipedia.org/wiki/Walter_Ulbricht
Walter van Tilburg Clark	http://en.wikipedia.org/wiki/Walter_van_Tilburg_Clark
Walter Wanger	http://en.wikipedia.org/wiki/Walter_Wanger
Walter Winchell	http://en.wikipedia.org/wiki/Walter_Winchell
Walther Bothe	http://en.wikipedia.org/wiki/Walther_Bothe
Walther Funk	http://en.wikipedia.org/wiki/Walther_Funk
Walther Nernst	http://en.wikipedia.org/wiki/Walther_Nernst
Walther von Brauchitsch	http://en.wikipedia.org/wiki/Walther_von_Brauchitsch
Walther von der Vogelweide	http://en.wikipedia.org/wiki/Walther_von_der_Vogelweide
Walther von Reichenau	http://en.wikipedia.org/wiki/Walther_von_Reichenau
Wanda Hendrix	http://en.wikipedia.org/wiki/Wanda_Hendrix
Wanda Sykes	http://en.wikipedia.org/wiki/Wanda_Sykes
Wang An	http://en.wikipedia.org/wiki/Wang_An
Wangari Maathai	http://en.wikipedia.org/wiki/Wangari_Maathai
Ward Bond	http://en.wikipedia.org/wiki/Ward_Bond
Ward Churchill	http://en.wikipedia.org/wiki/Ward_Churchill
Wardell Gray	http://en.wikipedia.org/wiki/Wardell_Gray
Warner Baxter	http://en.wikipedia.org/wiki/Warner_Baxter
Warner Oland	http://en.wikipedia.org/wiki/Warner_Oland
Warren B. Rudman	http://en.wikipedia.org/wiki/Warren_B._Rudman
Warren Barker	http://en.wikipedia.org/wiki/Warren_Barker
Warren Beatty	http://en.wikipedia.org/wiki/Warren_Beatty
Warren Bennis	http://en.wikipedia.org/wiki/Warren_Bennis
Warren Buffett	http://en.wikipedia.org/wiki/Warren_Buffett
Warren Burger	http://en.wikipedia.org/wiki/Warren_Burger
Warren Christopher	http://en.wikipedia.org/wiki/Warren_Christopher
Warren Ellis	http://en.wikipedia.org/wiki/Warren_Ellis
Warren G	http://en.wikipedia.org/wiki/Warren_G
Warren G. Harding	http://en.wikipedia.org/wiki/Warren_G._Harding
Warren Hastings	http://en.wikipedia.org/wiki/Warren_Hastings
Warren Hinckle	http://en.wikipedia.org/wiki/Warren_Hinckle
Warren Jeffs	http://en.wikipedia.org/wiki/Warren_Jeffs
Warren Oates	http://en.wikipedia.org/wiki/Warren_Oates
Warren Olney	http://en.wikipedia.org/wiki/Warren_Olney_(journalist)
Warren R. Austin	http://en.wikipedia.org/wiki/Warren_R._Austin
Warren Robinett	http://en.wikipedia.org/wiki/Warren_Robinett
Warren Rudman	http://en.wikipedia.org/wiki/Warren_Rudman
Warren Spahn	http://en.wikipedia.org/wiki/Warren_Spahn
Warren Zevon	http://en.wikipedia.org/wiki/Warren_Zevon
Warwick Davis	http://en.wikipedia.org/wiki/Warwick_Davis
Washington Allston	http://en.wikipedia.org/wiki/Washington_Allston
Washington Irving	http://en.wikipedia.org/wiki/Washington_Irving
Wassily Kandinsky	http://en.wikipedia.org/wiki/Wassily_Kandinsky
Wassily Leontief	http://en.wikipedia.org/wiki/Wassily_Leontief
Wat Tyler	http://en.wikipedia.org/wiki/Wat_Tyler
Wavy Gravy	http://en.wikipedia.org/wiki/Wavy_Gravy
Waylon Jennings	http://en.wikipedia.org/wiki/Waylon_Jennings
Wayne Allard	http://en.wikipedia.org/wiki/Wayne_Allard
Wayne Allyn Root	http://en.wikipedia.org/wiki/Wayne_Allyn_Root
Wayne Brady	http://en.wikipedia.org/wiki/Wayne_Brady
Wayne C. Booth	http://en.wikipedia.org/wiki/Wayne_C._Booth
Wayne Coyne	http://en.wikipedia.org/wiki/Wayne_Coyne
Wayne David	http://en.wikipedia.org/wiki/Wayne_David
Wayne Dowdy	http://en.wikipedia.org/wiki/Wayne_Dowdy
Wayne Dyer	http://en.wikipedia.org/wiki/Wayne_Dyer
Wayne Gilchrest	http://en.wikipedia.org/wiki/Wayne_Gilchrest
Wayne Gretzky	http://en.wikipedia.org/wiki/Wayne_Gretzky
Wayne Knight	http://en.wikipedia.org/wiki/Wayne_Knight
Wayne LaPierre	http://en.wikipedia.org/wiki/Wayne_LaPierre
Wayne Newton	http://en.wikipedia.org/wiki/Wayne_Newton
Wayne Osmond	http://en.wikipedia.org/wiki/Wayne_Osmond
Wayne Rogers	http://en.wikipedia.org/wiki/Wayne_Rogers
Wayne Rooney	http://en.wikipedia.org/wiki/Wayne_Rooney
Wayne Thiebaud	http://en.wikipedia.org/wiki/Wayne_Thiebaud
Wayne Wang	http://en.wikipedia.org/wiki/Wayne_Wang
Wayne Williams	http://en.wikipedia.org/wiki/Wayne_Williams
Wayne Wonder	http://en.wikipedia.org/wiki/Wayne_Wonder
Webb Franklin	http://en.wikipedia.org/wiki/Webb_Franklin
Webb Hubbell	http://en.wikipedia.org/wiki/Webb_Hubbell
Weird Al Yankovic	http://en.wikipedia.org/wiki/Weird_Al_Yankovic
Wellington Mara	http://en.wikipedia.org/wiki/Wellington_Mara
Wen Ho Lee	http://en.wikipedia.org/wiki/Wen_Ho_Lee
Wen Jiabao	http://en.wikipedia.org/wiki/Wen_Jiabao
Wendell Berry	http://en.wikipedia.org/wiki/Wendell_Berry
Wendell Corey	http://en.wikipedia.org/wiki/Wendell_Corey
Wendell H. Ford	http://en.wikipedia.org/wiki/Wendell_H._Ford
Wendell M. Stanley	http://en.wikipedia.org/wiki/Wendell_M._Stanley
Wendell Willkie	http://en.wikipedia.org/wiki/Wendell_Willkie
Wendi McLendon-Covey	http://en.wikipedia.org/wiki/Wendi_McLendon-Covey
Wendie Jo Sperber	http://en.wikipedia.org/wiki/Wendie_Jo_Sperber
Wendie Malick	http://en.wikipedia.org/wiki/Wendie_Malick
Wendy Carlos	http://en.wikipedia.org/wiki/Wendy_Carlos
Wendy Cope	http://en.wikipedia.org/wiki/Wendy_Cope
Wendy Crewson	http://en.wikipedia.org/wiki/Wendy_Crewson
Wendy Gramm	http://en.wikipedia.org/wiki/Wendy_Gramm
Wendy Hiller	http://en.wikipedia.org/wiki/Wendy_Hiller
Wendy Makkena	http://en.wikipedia.org/wiki/Wendy_Makkena
Wendy O. Williams	http://en.wikipedia.org/wiki/Wendy_O._Williams
Wendy Pini	http://en.wikipedia.org/wiki/Wendy_Pini
Wendy Wasserstein	http://en.wikipedia.org/wiki/Wendy_Wasserstein
Wentworth Miller	http://en.wikipedia.org/wiki/Wentworth_Miller
Wenzel Hollar	http://en.wikipedia.org/wiki/Wenzel_Hollar
Werner Erhard	http://en.wikipedia.org/wiki/Werner_Erhard
Werner Faymann	http://en.wikipedia.org/wiki/Werner_Faymann
Werner Heisenberg	http://en.wikipedia.org/wiki/Werner_Heisenberg
Werner Herzog	http://en.wikipedia.org/wiki/Werner_Herzog
Werner Klemperer	http://en.wikipedia.org/wiki/Werner_Klemperer
Werner von Blomberg	http://en.wikipedia.org/wiki/Werner_von_Blomberg
Wernher von Braun	http://en.wikipedia.org/wiki/Wernher_von_Braun
Wes Anderson	http://en.wikipedia.org/wiki/Wes_Anderson
Wes Bentley	http://en.wikipedia.org/wiki/Wes_Bentley
Wes Boyd	http://en.wikipedia.org/wiki/Wes_Boyd
Wes Craven	http://en.wikipedia.org/wiki/Wes_Craven
Wes Montgomery	http://en.wikipedia.org/wiki/Wes_Montgomery
Wes Pruden	http://en.wikipedia.org/wiki/Wes_Pruden
Wes Studi	http://en.wikipedia.org/wiki/Wes_Studi
Wes Watkins	http://en.wikipedia.org/wiki/Wes_Watkins
Wesley Addy	http://en.wikipedia.org/wiki/Wesley_Addy
Wesley Clark	http://en.wikipedia.org/wiki/Wesley_Clark
Wesley Snipes	http://en.wikipedia.org/wiki/Wesley_Snipes
Wesley Willis	http://en.wikipedia.org/wiki/Wesley_Willis
Whit Bissell	http://en.wikipedia.org/wiki/Whit_Bissell
Whitey Bulger	http://en.wikipedia.org/wiki/Whitey_Bulger
Whitey Ford	http://en.wikipedia.org/wiki/Whitey_Ford
Whitey Herzog	http://en.wikipedia.org/wiki/Whitey_Herzog
Whitfield Diffie	http://en.wikipedia.org/wiki/Whitfield_Diffie
Whitley Strieber	http://en.wikipedia.org/wiki/Whitley_Strieber
Whitney Houston	http://en.wikipedia.org/wiki/Whitney_Houston
Whittaker Chambers	http://en.wikipedia.org/wiki/Whittaker_Chambers
Whoopi Goldberg	http://en.wikipedia.org/wiki/Whoopi_Goldberg
Wietse Venema	http://en.wikipedia.org/wiki/Wietse_Venema
Wil Wheaton	http://en.wikipedia.org/wiki/Wil_Wheaton
Wilbert Harrison	http://en.wikipedia.org/wiki/Wilbert_Harrison
Wilbert J. "Billy" Tauzin	http://en.wikipedia.org/wiki/Wilbert_J._%22Billy%22_Tauzin
Wilbur Ross	http://en.wikipedia.org/wiki/Wilbur_Ross
Wilbur Scoville	http://en.wikipedia.org/wiki/Wilbur_Scoville
Wilbur Wright	http://en.wikipedia.org/wiki/Wilbur_Wright
Wild Bill Donovan	http://en.wikipedia.org/wiki/Wild_Bill_Donovan
Wild Bill Elliott	http://en.wikipedia.org/wiki/Wild_Bill_Elliott
Wild Bill Hickok	http://en.wikipedia.org/wiki/Wild_Bill_Hickok
Wilds Preston Richardson	http://en.wikipedia.org/wiki/Wilds_Preston_Richardson
Wiley Post	http://en.wikipedia.org/wiki/Wiley_Post
Wilford B. Hoggatt	http://en.wikipedia.org/wiki/Wilford_B._Hoggatt
Wilford Brimley	http://en.wikipedia.org/wiki/Wilford_Brimley
Wilfred Owen	http://en.wikipedia.org/wiki/Wilfred_Owen
Wilfrid Laurier	http://en.wikipedia.org/wiki/Wilfrid_Laurier
Wilfrid Sheed	http://en.wikipedia.org/wiki/Wilfrid_Sheed
Wilhelm Canaris	http://en.wikipedia.org/wiki/Wilhelm_Canaris
Wilhelm Conrad R�ntgen	http://en.wikipedia.org/wiki/Wilhelm_Conrad_R%F6ntgen
Wilhelm Cuno	http://en.wikipedia.org/wiki/Wilhelm_Cuno
Wilhelm Frick	http://en.wikipedia.org/wiki/Wilhelm_Frick
Wilhelm Furtw�ngler	http://en.wikipedia.org/wiki/Wilhelm_Furtw%E4ngler
Wilhelm Hauff	http://en.wikipedia.org/wiki/Wilhelm_Hauff
Wilhelm Hofmeister	http://en.wikipedia.org/wiki/Wilhelm_Hofmeister
Wilhelm Junker	http://en.wikipedia.org/wiki/Wilhelm_Junker
Wilhelm Keitel	http://en.wikipedia.org/wiki/Wilhelm_Keitel
Wilhelm Marx	http://en.wikipedia.org/wiki/Wilhelm_Marx
Wilhelm Olbers	http://en.wikipedia.org/wiki/Wilhelm_Olbers
Wilhelm Ostwald	http://en.wikipedia.org/wiki/Wilhelm_Ostwald
Wilhelm Pieck	http://en.wikipedia.org/wiki/Wilhelm_Pieck
Wilhelm Reich	http://en.wikipedia.org/wiki/Wilhelm_Reich
Wilhelm von Humboldt	http://en.wikipedia.org/wiki/Wilhelm_von_Humboldt
Wilhelm Weber	http://en.wikipedia.org/wiki/Wilhelm_Eduard_Weber
Wilhelm Wien	http://en.wikipedia.org/wiki/Wilhelm_Wien
Wilhelm Wundt	http://en.wikipedia.org/wiki/Wilhelm_Wundt
Wilkie Collins	http://en.wikipedia.org/wiki/Wilkie_Collins
Will Arnett	http://en.wikipedia.org/wiki/Will_Arnett
Will Durant	http://en.wikipedia.org/wiki/Will_Durant
Will Eisner	http://en.wikipedia.org/wiki/Will_Eisner
Will Estes	http://en.wikipedia.org/wiki/Will_Estes
Will Ferrell	http://en.wikipedia.org/wiki/Will_Ferrell
Will Forte	http://en.wikipedia.org/wiki/Will_Forte
Will Friedle	http://en.wikipedia.org/wiki/Will_Friedle
Will Geer	http://en.wikipedia.org/wiki/Will_Geer
Will Hay	http://en.wikipedia.org/wiki/Will_Hay
Will Hutchins	http://en.wikipedia.org/wiki/Will_Hutchins
Will Oldham	http://en.wikipedia.org/wiki/Will_Oldham
Will Patton	http://en.wikipedia.org/wiki/Will_Patton
Will Rogers	http://en.wikipedia.org/wiki/Will_Rogers
Will Rogers, Jr.	http://en.wikipedia.org/wiki/Will_Rogers%2C_Jr.
Will Rothhaar	http://en.wikipedia.org/wiki/Will_Rothhaar
Will Sasso	http://en.wikipedia.org/wiki/Will_Sasso
Will Sergeant	http://en.wikipedia.org/wiki/Will_Sergeant
Will Smith	http://en.wikipedia.org/wiki/Will_Smith
Will Wright	http://en.wikipedia.org/wiki/Will_Wright_(game_designer)
Will Young	http://en.wikipedia.org/wiki/Will_Young
Willa Cather	http://en.wikipedia.org/wiki/Willa_Cather
Willard F. Libby	http://en.wikipedia.org/wiki/Willard_F._Libby
Willard Scott	http://en.wikipedia.org/wiki/Willard_Scott
Willard Van Orman Quine	http://en.wikipedia.org/wiki/Willard_Van_Orman_Quine
Willard Wirtz	http://en.wikipedia.org/wiki/Willard_Wirtz
Willem Barents	http://en.wikipedia.org/wiki/Willem_Barents
Willem Dafoe	http://en.wikipedia.org/wiki/Willem_Dafoe
Willem de Kooning	http://en.wikipedia.org/wiki/Willem_de_Kooning
Willi Stoph	http://en.wikipedia.org/wiki/Willi_Stoph
William "The Refrigerator" Perry	http://en.wikipedia.org/wiki/William_%22The_Refrigerator%22_Perry
William A. Fowler	http://en.wikipedia.org/wiki/William_A._Fowler
William A. O'Neill	http://en.wikipedia.org/wiki/William_A._O%27Neill
William A. Osborn	http://en.wikipedia.org/wiki/William_A._Osborn
William A. Seiter	http://en.wikipedia.org/wiki/William_A._Seiter
William A. Wellman	http://en.wikipedia.org/wiki/William_A._Wellman
William A. Wheeler	http://en.wikipedia.org/wiki/William_A._Wheeler
William Allen White	http://en.wikipedia.org/wiki/William_Allen_White
William Allingham	http://en.wikipedia.org/wiki/William_Allingham
William Apess	http://en.wikipedia.org/wiki/William_Apess
William B. Davis	http://en.wikipedia.org/wiki/William_B._Davis
William B. Harrison Jr.	http://en.wikipedia.org/wiki/William_B._Harrison,_Jr.
William Baffin	http://en.wikipedia.org/wiki/William_Baffin
William Bagley	http://en.wikipedia.org/wiki/William_Bagley_(educator)
William Bain	http://en.wikipedia.org/wiki/Willie_Bain
William Bainbridge	http://en.wikipedia.org/wiki/William_Bainbridge
William Baldwin	http://en.wikipedia.org/wiki/William_Baldwin
William Barker Cushing	http://en.wikipedia.org/wiki/William_Barker_Cushing
William Barr	http://en.wikipedia.org/wiki/William_Barr_(politician)
William Bartram	http://en.wikipedia.org/wiki/William_Bartram
William Bateson	http://en.wikipedia.org/wiki/William_Bateson
William Bayliss	http://en.wikipedia.org/wiki/William_Bayliss
William Bendix	http://en.wikipedia.org/wiki/William_Bendix
William Bennett	http://en.wikipedia.org/wiki/William_Bennett
William Bennett	http://en.wikipedia.org/wiki/William_Bennett
William Blackstone	http://en.wikipedia.org/wiki/William_Blackstone
William Blake	http://en.wikipedia.org/wiki/William_Blake
William Booth	http://en.wikipedia.org/wiki/William_Booth
William Boyce	http://en.wikipedia.org/wiki/William_Boyce
William Boyd	http://en.wikipedia.org/wiki/William_Boyd_(actor)
William Boyd Allison	http://en.wikipedia.org/wiki/William_Boyd_Allison
William Bradford	http://en.wikipedia.org/wiki/William_Bradford_(Colonial_printer)
William Bradford	http://en.wikipedia.org/wiki/William_Bradford_(Plymouth_governor)
William Bragg	http://en.wikipedia.org/wiki/William_Henry_Bragg
William Brockman Bankhead	http://en.wikipedia.org/wiki/William_Brockman_Bankhead
William Buckland	http://en.wikipedia.org/wiki/William_Buckland
William Bulow	http://en.wikipedia.org/wiki/William_Bulow
William Bundy	http://en.wikipedia.org/wiki/William_Bundy
William Burke	http://en.wikipedia.org/wiki/William_Burke
William Butler Yeats	http://en.wikipedia.org/wiki/William_Butler_Yeats
William Byrd	http://en.wikipedia.org/wiki/William_Byrd
William C. Bouck	http://en.wikipedia.org/wiki/William_C._Bouck
William C. Durant	http://en.wikipedia.org/wiki/William_C._Durant
William C. Weldon	http://en.wikipedia.org/wiki/William_C._Weldon
William C. Whitney	http://en.wikipedia.org/wiki/William_C._Whitney
William Calley	http://en.wikipedia.org/wiki/William_Calley
William Camden	http://en.wikipedia.org/wiki/William_Camden
William Carey	http://en.wikipedia.org/wiki/William_Carey_(missionary)
William Carlos Williams	http://en.wikipedia.org/wiki/William_Carlos_Williams
William Carney	http://en.wikipedia.org/wiki/William_Carney_(politician)
William Casey	http://en.wikipedia.org/wiki/William_Casey
William Cash	http://en.wikipedia.org/wiki/William_Cash
William Caslon	http://en.wikipedia.org/wiki/William_Caslon
William Castle	http://en.wikipedia.org/wiki/William_Castle
William Caxton	http://en.wikipedia.org/wiki/William_Caxton
William Cecil	http://en.wikipedia.org/wiki/William_Cecil,_1st_Baron_Burghley
William Chambers	http://en.wikipedia.org/wiki/William_Chambers_(publisher)
William Charles Macready	http://en.wikipedia.org/wiki/William_Charles_Macready
William Christopher	http://en.wikipedia.org/wiki/William_Christopher
William Clark	http://en.wikipedia.org/wiki/William_Clark_(explorer)
William Clay Ford, Jr.	http://en.wikipedia.org/wiki/William_Clay_Ford%2C_Jr.
William Clay Ford, Sr.	http://en.wikipedia.org/wiki/William_Clay_Ford%2C_Sr.
William Cobbett	http://en.wikipedia.org/wiki/William_Cobbett
William Cohen	http://en.wikipedia.org/wiki/William_Cohen
William Colby	http://en.wikipedia.org/wiki/William_Colby
William Congreve	http://en.wikipedia.org/wiki/William_Congreve
William Conrad	http://en.wikipedia.org/wiki/William_Conrad
William Cowper	http://en.wikipedia.org/wiki/William_Cowper
William Cullen Bryant	http://en.wikipedia.org/wiki/William_Cullen_Bryant
William D. Ford	http://en.wikipedia.org/wiki/William_D._Ford
William D. Ford	http://en.wikipedia.org/wiki/William_D._Ford
William D. Lutz	http://en.wikipedia.org/wiki/William_D._Lutz
William D. Phillips	http://en.wikipedia.org/wiki/William_D._Phillips
William Dampier	http://en.wikipedia.org/wiki/William_Dampier
William Daniels	http://en.wikipedia.org/wiki/William_Daniels
William Davison	http://en.wikipedia.org/wiki/William_Davison_(diplomat)
William Dean Howells	http://en.wikipedia.org/wiki/William_Dean_Howells
William Demarest	http://en.wikipedia.org/wiki/William_Demarest
William Desmond Taylor	http://en.wikipedia.org/wiki/William_Desmond_Taylor
William Devane	http://en.wikipedia.org/wiki/William_Devane
William Dieterle	http://en.wikipedia.org/wiki/William_Dieterle
William Dodd Hathaway	http://en.wikipedia.org/wiki/William_Dodd_Hathaway
William Donald Schaefer	http://en.wikipedia.org/wiki/William_Donald_Schaefer
William Donohue	http://en.wikipedia.org/wiki/William_Donohue
William Dunbar	http://en.wikipedia.org/wiki/William_Dunbar
William Dunlap	http://en.wikipedia.org/wiki/William_Dunlap
William E. Brock	http://en.wikipedia.org/wiki/William_E._Brock
William E. Dannemeyer	http://en.wikipedia.org/wiki/William_E._Dannemeyer
William E. Kennard	http://en.wikipedia.org/wiki/William_E._Kennard
William Edward Forster	http://en.wikipedia.org/wiki/William_Edward_Forster
William Empson	http://en.wikipedia.org/wiki/William_Empson
William Evans Burton	http://en.wikipedia.org/wiki/William_Evans_Burton
William Ewart Gladstone	http://en.wikipedia.org/wiki/William_Ewart_Gladstone
William F. Buckley	http://en.wikipedia.org/wiki/William_F._Buckley
William F. Clinger	http://en.wikipedia.org/wiki/William_F._Clinger
William F. Giauque	http://en.wikipedia.org/wiki/William_F._Giauque
William F. Goodling	http://en.wikipedia.org/wiki/William_F._Goodling
William F. Halsey	http://en.wikipedia.org/wiki/William_F._Halsey
William F. Harrah	http://en.wikipedia.org/wiki/William_F._Harrah
William F. Raborn	http://en.wikipedia.org/wiki/William_Raborn
William Faulkner	http://en.wikipedia.org/wiki/William_Faulkner
William Forsythe	http://en.wikipedia.org/wiki/William_Forsythe_(actor)
William Foxwell Albright	http://en.wikipedia.org/wiki/William_Foxwell_Albright
William Frawley	http://en.wikipedia.org/wiki/William_Frawley
William French Smith	http://en.wikipedia.org/wiki/William_French_Smith
William Friedkin	http://en.wikipedia.org/wiki/William_Friedkin
William Friedman	http://en.wikipedia.org/wiki/William_Friedman
William Gaddis	http://en.wikipedia.org/wiki/William_Gaddis
William Gibson	http://en.wikipedia.org/wiki/William_Gibson
William Gilbert	http://en.wikipedia.org/wiki/William_Gilbert
William Gillette	http://en.wikipedia.org/wiki/William_Gillette
William Godwin	http://en.wikipedia.org/wiki/William_Godwin
William Golding	http://en.wikipedia.org/wiki/William_Golding
William Goldman	http://en.wikipedia.org/wiki/William_Goldman
William Goldman	http://en.wikipedia.org/wiki/William_Goldman
William Grayson	http://en.wikipedia.org/wiki/William_Grayson
William H. Crawford	http://en.wikipedia.org/wiki/William_H._Crawford
William H. Gass	http://en.wikipedia.org/wiki/William_H._Gass
William H. Gray	http://en.wikipedia.org/wiki/William_H._Gray_(congressman)
William H. Gray, III	http://en.wikipedia.org/wiki/William_H._Gray_(congressman)
William H. Macy	http://en.wikipedia.org/wiki/William_H._Macy
William H. Natcher	http://en.wikipedia.org/wiki/William_H._Natcher
William H. Natcher	http://en.wikipedia.org/wiki/William_H._Natcher
William H. Stein	http://en.wikipedia.org/wiki/William_H._Stein
William Habington	http://en.wikipedia.org/wiki/William_Habington
William Hague	http://en.wikipedia.org/wiki/William_Hague
William Haines	http://en.wikipedia.org/wiki/William_Haines
William Hanna	http://en.wikipedia.org/wiki/William_Hanna
William Harrison	http://en.wikipedia.org/wiki/William_B._Harrison,_Jr.
William Harrison Ainsworth	http://en.wikipedia.org/wiki/William_Harrison_Ainsworth
William Hartnell	http://en.wikipedia.org/wiki/William_Hartnell
William Harvey	http://en.wikipedia.org/wiki/William_Harvey
William Hazlitt	http://en.wikipedia.org/wiki/William_Hazlitt
William Henry	http://en.wikipedia.org/wiki/William_Henry_(chemist)
William Henry Ashley	http://en.wikipedia.org/wiki/William_Henry_Ashley
William Henry Davies	http://en.wikipedia.org/wiki/William_Henry_Davies
William Henry Fox Talbot	http://en.wikipedia.org/wiki/William_Henry_Fox_Talbot
William Henry Harrison	http://en.wikipedia.org/wiki/William_Henry_Harrison
William Henry Ireland	http://en.wikipedia.org/wiki/William_Henry_Ireland
William Henry Perkin	http://en.wikipedia.org/wiki/William_Henry_Perkin
William Henry Seward	http://en.wikipedia.org/wiki/William_Henry_Seward
William Henry Vanderbilt	http://en.wikipedia.org/wiki/William_Henry_Vanderbilt
William Herschel	http://en.wikipedia.org/wiki/William_Herschel
William Hewlett	http://en.wikipedia.org/wiki/William_Reddington_Hewlett
William Hogarth	http://en.wikipedia.org/wiki/William_Hogarth
William Holden	http://en.wikipedia.org/wiki/William_Holden
William Holman Hunt	http://en.wikipedia.org/wiki/William_Holman_Hunt
William Hone	http://en.wikipedia.org/wiki/William_Hone
William Hopper	http://en.wikipedia.org/wiki/William_Hopper
William Horsley	http://en.wikipedia.org/wiki/William_Horsley
William Hoste	http://en.wikipedia.org/wiki/William_Hoste
William Hotham	http://en.wikipedia.org/wiki/William_Hotham_(1772_-_1848)
William Howard Taft	http://en.wikipedia.org/wiki/William_Howard_Taft
William Howe	http://en.wikipedia.org/wiki/William_Howe,_5th_Viscount_Howe
William Howitt	http://en.wikipedia.org/wiki/William_Howitt
William Huggins	http://en.wikipedia.org/wiki/William_Huggins
William Hung	http://en.wikipedia.org/wiki/William_Hung
William Hunter	http://en.wikipedia.org/wiki/William_Hunter_(anatomist)
William Hurt	http://en.wikipedia.org/wiki/William_Hurt
William Hyde Wollaston	http://en.wikipedia.org/wiki/William_Hyde_Wollaston
William Inge	http://en.wikipedia.org/wiki/William_Inge
William J. B. Dorn	http://en.wikipedia.org/wiki/William_Jennings_Bryan_Dorn
William J. Brennan	http://en.wikipedia.org/wiki/William_J._Brennan
William J. Burns	http://en.wikipedia.org/wiki/William_J._Burns
William J. Coyne	http://en.wikipedia.org/wiki/William_J._Coyne
William J. Flynn	http://en.wikipedia.org/wiki/William_J._Flynn
William J. Hughes	http://en.wikipedia.org/wiki/William_J._Hughes
William J. Lynn III	http://en.wikipedia.org/wiki/William_J._Lynn_III
William J. Perry	http://en.wikipedia.org/wiki/William_J._Perry
William Jackson Hooker	http://en.wikipedia.org/wiki/William_Jackson_Hooker
William James	http://en.wikipedia.org/wiki/William_James
William James Mayo	http://en.wikipedia.org/wiki/William_James_Mayo
William Jefferson	http://en.wikipedia.org/wiki/William_J._Jefferson
William Jennings Bryan	http://en.wikipedia.org/wiki/William_Jennings_Bryan
William Joseph Hardee	http://en.wikipedia.org/wiki/William_Joseph_Hardee
William Julius Wilson	http://en.wikipedia.org/wiki/William_Julius_Wilson
William Katt	http://en.wikipedia.org/wiki/William_Katt
William Keighley	http://en.wikipedia.org/wiki/William_Keighley
William Kennedy	http://en.wikipedia.org/wiki/William_Joseph_Kennedy
William Kennedy Smith	http://en.wikipedia.org/wiki/William_Kennedy_Smith
William Kent	http://en.wikipedia.org/wiki/William_Kent
William Kunstler	http://en.wikipedia.org/wiki/William_Kunstler
William L. Armstrong	http://en.wikipedia.org/wiki/William_L._Armstrong
William L. Clay	http://en.wikipedia.org/wiki/William_L._Clay
William L. Clay	http://en.wikipedia.org/wiki/William_L._Clay
William L. Marcy	http://en.wikipedia.org/wiki/William_L._Marcy
William L. Petersen	http://en.wikipedia.org/wiki/William_L._Petersen
William L. Shirer	http://en.wikipedia.org/wiki/William_L._Shirer
William Langer	http://en.wikipedia.org/wiki/William_Langer
William Laud	http://en.wikipedia.org/wiki/William_Laud
William Law	http://en.wikipedia.org/wiki/William_Law
William Lawrence Allen	http://en.wikipedia.org/wiki/William_Lawrence_Allen
William Least Heat-Moon	http://en.wikipedia.org/wiki/William_Least_Heat-Moon
William Lehman	http://en.wikipedia.org/wiki/William_Lehman_(Florida_politician)
William Leonard	http://en.wikipedia.org/wiki/William_J._Leonard
William Leonard Langer	http://en.wikipedia.org/wiki/William_Leonard_Langer
William Levitt	http://en.wikipedia.org/wiki/William_Levitt
William Lipscomb	http://en.wikipedia.org/wiki/William_Lipscomb
William Lloyd Garrison	http://en.wikipedia.org/wiki/William_Lloyd_Garrison
William Lundigan	http://en.wikipedia.org/wiki/William_Lundigan
William Lyon Mackenzie King	http://en.wikipedia.org/wiki/William_Lyon_Mackenzie_King
William Lyon Phelps	http://en.wikipedia.org/wiki/William_Lyon_Phelps
William M. Daley	http://en.wikipedia.org/wiki/William_M._Daley
William M. Evarts	http://en.wikipedia.org/wiki/William_M._Evarts
William Makepeace Thackeray	http://en.wikipedia.org/wiki/William_Makepeace_Thackeray
William Manchester	http://en.wikipedia.org/wiki/William_Manchester
William Mapother	http://en.wikipedia.org/wiki/William_Mapother
William Marshall	http://en.wikipedia.org/wiki/William_Marshall_(bandleader)
William Masters	http://en.wikipedia.org/wiki/William_Masters
William Maxwell	http://en.wikipedia.org/wiki/William_Keepers_Maxwell,_Jr.
William McChesney Martin	http://en.wikipedia.org/wiki/William_McChesney_Martin
William McCrea	http://en.wikipedia.org/wiki/William_McCrea_(politician)
William McDonough	http://en.wikipedia.org/wiki/William_McDonough
William McDougall	http://en.wikipedia.org/wiki/William_McDougall_(psychologist)
William McKinley	http://en.wikipedia.org/wiki/William_McKinley
William McNamara	http://en.wikipedia.org/wiki/William_McNamara
William Meredith	http://en.wikipedia.org/wiki/William_Morris_Meredith,_Jr.
William Monroe Trotter	http://en.wikipedia.org/wiki/William_Monroe_Trotter
William Moon	http://en.wikipedia.org/wiki/William_Moon
William Morris	http://en.wikipedia.org/wiki/William_Morris
William Morris	http://en.wikipedia.org/wiki/William_N._Morris
William Moseley	http://en.wikipedia.org/wiki/William_Moseley_(actor)
William Moulton Marston	http://en.wikipedia.org/wiki/William_Moulton_Marston
William Niskanen	http://en.wikipedia.org/wiki/William_Niskanen
William O. Douglas	http://en.wikipedia.org/wiki/William_O._Douglas
William O. Lipinski	http://en.wikipedia.org/wiki/William_O._Lipinski
William O. Studeman	http://en.wikipedia.org/wiki/William_O._Studeman
William Odom	http://en.wikipedia.org/wiki/William_Odom
William of Ockham	http://en.wikipedia.org/wiki/William_of_Ockham
William of Orange	http://en.wikipedia.org/wiki/William_III_of_England
William Osler	http://en.wikipedia.org/wiki/William_Osler
William Oughtred	http://en.wikipedia.org/wiki/William_Oughtred
William P. Clark	http://en.wikipedia.org/wiki/William_P._Clark
William P. Lauder	http://en.wikipedia.org/wiki/William_P._Lauder
William P. Lear	http://en.wikipedia.org/wiki/William_P._Lear
William P. Rogers	http://en.wikipedia.org/wiki/William_P._Rogers
William Paley	http://en.wikipedia.org/wiki/William_Paley
William Paterson	http://en.wikipedia.org/wiki/William_Paterson_(banker)
William Paterson	http://en.wikipedia.org/wiki/William_Paterson_(judge)
William Penn	http://en.wikipedia.org/wiki/William_Penn
William Peter Blatty	http://en.wikipedia.org/wiki/William_Peter_Blatty
William Pierce	http://en.wikipedia.org/wiki/William_Luther_Pierce
William Pitt the Younger	http://en.wikipedia.org/wiki/William_Pitt_the_Younger
William Powell	http://en.wikipedia.org/wiki/William_Powell
William Proxmire	http://en.wikipedia.org/wiki/William_Proxmire
William Proxmire	http://en.wikipedia.org/wiki/William_Proxmire
William R. King	http://en.wikipedia.org/wiki/William_R._King
William R. Moses	http://en.wikipedia.org/wiki/William_R._Moses
William Randolph Hearst	http://en.wikipedia.org/wiki/William_Randolph_Hearst
William Rehnquist	http://en.wikipedia.org/wiki/William_Rehnquist
William Robertson	http://en.wikipedia.org/wiki/William_Robertson
William Rose Ben�t	http://en.wikipedia.org/wiki/William_Rose_Ben%E9t
William Rosenberg	http://en.wikipedia.org/wiki/William_Rosenberg
William Rowley	http://en.wikipedia.org/wiki/William_Rowley
William Ruckelshaus	http://en.wikipedia.org/wiki/William_Ruckelshaus
William Russ	http://en.wikipedia.org/wiki/William_Russ
William Ryan	http://en.wikipedia.org/wiki/William_Ryan
William S. Broomfield	http://en.wikipedia.org/wiki/William_S._Broomfield
William S. Burroughs	http://en.wikipedia.org/wiki/William_S._Burroughs
William S. Cohen	http://en.wikipedia.org/wiki/William_S._Cohen
William S. Farish	http://en.wikipedia.org/wiki/William_Stamps_Farish_III
William S. Hart	http://en.wikipedia.org/wiki/William_S._Hart
William S. Knowles	http://en.wikipedia.org/wiki/William_S._Knowles
William S. Paley	http://en.wikipedia.org/wiki/William_S._Paley
William S. Rosecrans	http://en.wikipedia.org/wiki/William_S._Rosecrans
William S. Rukeyser	http://en.wikipedia.org/wiki/William_S._Rukeyser
William Safire	http://en.wikipedia.org/wiki/William_Safire
William Sanderson	http://en.wikipedia.org/wiki/William_Sanderson
William Saroyan	http://en.wikipedia.org/wiki/William_Saroyan
William Schreyer	http://en.wikipedia.org/wiki/William_Schreyer
William Schuman	http://en.wikipedia.org/wiki/William_Schuman
William Seabrook	http://en.wikipedia.org/wiki/William_Seabrook
William Sessions	http://en.wikipedia.org/wiki/William_S._Sessions
William Shakespeare	http://en.wikipedia.org/wiki/William_Shakespeare
William Shatner	http://en.wikipedia.org/wiki/William_Shatner
William Shawn	http://en.wikipedia.org/wiki/William_Shawn
William Shenstone	http://en.wikipedia.org/wiki/William_Shenstone
William Shirley	http://en.wikipedia.org/wiki/William_Shirley
William Shockley	http://en.wikipedia.org/wiki/William_Shockley
William Sloane Coffin	http://en.wikipedia.org/wiki/William_Sloane_Coffin
William Smith	http://en.wikipedia.org/wiki/William_Smith_(geologist)
William Snow Harris	http://en.wikipedia.org/wiki/William_Snow_Harris
William Stafford	http://en.wikipedia.org/wiki/William_Stafford_(poet)
William Stanley Jevons	http://en.wikipedia.org/wiki/William_Stanley_Jevons
William Steig	http://en.wikipedia.org/wiki/William_Steig
William Strode	http://en.wikipedia.org/wiki/William_Strode
William Stubbs	http://en.wikipedia.org/wiki/William_Stubbs
William Stukeley	http://en.wikipedia.org/wiki/William_Stukeley
William Styron	http://en.wikipedia.org/wiki/William_Styron
William T. Orr	http://en.wikipedia.org/wiki/William_T._Orr
William T. Sherman	http://en.wikipedia.org/wiki/William_T._Sherman
William T. Vollmann	http://en.wikipedia.org/wiki/William_T._Vollmann
William Taylor Adams	http://en.wikipedia.org/wiki/William_Taylor_Adams
William the Conqueror	http://en.wikipedia.org/wiki/William_the_Conqueror
William Thomas Beckford	http://en.wikipedia.org/wiki/William_Thomas_Beckford
William Torrey Harris	http://en.wikipedia.org/wiki/William_Torrey_Harris
William Trevor	http://en.wikipedia.org/wiki/William_Trevor
William Trotter Bush	http://en.wikipedia.org/wiki/William_H._T._Bush
William Tyndale	http://en.wikipedia.org/wiki/William_Tyndale
William V. Roth, Jr.	http://en.wikipedia.org/wiki/William_V._Roth%2C_Jr.
William Vaughn Moody	http://en.wikipedia.org/wiki/William_Vaughn_Moody
William Walker	http://en.wikipedia.org/wiki/William_Walker_(filibuster)
William Wallace	http://en.wikipedia.org/wiki/William_Wallace
William Walsh	http://en.wikipedia.org/wiki/William_Walsh_(poet)
William Walton	http://en.wikipedia.org/wiki/William_Walton
William Warburton	http://en.wikipedia.org/wiki/William_Warburton
William Warham	http://en.wikipedia.org/wiki/William_Warham
William Weaver	http://en.wikipedia.org/wiki/William_Weaver
William Webster	http://en.wikipedia.org/wiki/William_H._Webster
William Westmoreland	http://en.wikipedia.org/wiki/William_Westmoreland
William Wetmore Story	http://en.wikipedia.org/wiki/William_Wetmore_Story
William Wharton	http://en.wikipedia.org/wiki/William_Wharton_(author)
William Whiston	http://en.wikipedia.org/wiki/William_Whiston
William Wilberforce	http://en.wikipedia.org/wiki/William_Wilberforce
William Windom	http://en.wikipedia.org/wiki/William_Windom
William Wirt	http://en.wikipedia.org/wiki/William_Wirt_(Attorney_General)
William Wollaston	http://en.wikipedia.org/wiki/William_Wollaston
William Wordsworth	http://en.wikipedia.org/wiki/William_Wordsworth
William Wycherley	http://en.wikipedia.org/wiki/William_Wycherley
William Wyler	http://en.wikipedia.org/wiki/William_Wyler
William Wyndham Grenville	http://en.wikipedia.org/wiki/William_Wyndham_Grenville
Willie Aames	http://en.wikipedia.org/wiki/Willie_Aames
Willie Bosket	http://en.wikipedia.org/wiki/Willie_Bosket
Willie Brown	http://en.wikipedia.org/wiki/Willie_Brown_(politician)
Willie D. Davis	http://en.wikipedia.org/wiki/Willie_Davis_(defensive_end)
Willie Garson	http://en.wikipedia.org/wiki/Willie_Garson
Willie Herenton	http://en.wikipedia.org/wiki/Willie_Herenton
Willie Horton	http://en.wikipedia.org/wiki/Willie_Horton
Willie Mays	http://en.wikipedia.org/wiki/Willie_Mays
Willie McCovey	http://en.wikipedia.org/wiki/Willie_McCovey
Willie Morris	http://en.wikipedia.org/wiki/Willie_Morris
Willie Mosconi	http://en.wikipedia.org/wiki/Willie_Mosconi
Willie Nelson	http://en.wikipedia.org/wiki/Willie_Nelson
Willie Shoemaker	http://en.wikipedia.org/wiki/Willie_Shoemaker
Willie Stargell	http://en.wikipedia.org/wiki/Willie_Stargell
Willie Sutton	http://en.wikipedia.org/wiki/Willie_Sutton
Willie Tyler	http://en.wikipedia.org/wiki/Willie_Tyler
Willis Carrier	http://en.wikipedia.org/wiki/Willis_Carrier
Willis D. Gradison Jr.	http://en.wikipedia.org/wiki/Willis_D._Gradison_Jr.
Willis Lamb	http://en.wikipedia.org/wiki/Willis_Lamb
Willy Brandt	http://en.wikipedia.org/wiki/Willy_Brandt
Willy Ley	http://en.wikipedia.org/wiki/Willy_Ley
Wilma Rudolph	http://en.wikipedia.org/wiki/Wilma_Rudolph
Wilmer Valderrama	http://en.wikipedia.org/wiki/Wilmer_Valderrama
Wilson Harris	http://en.wikipedia.org/wiki/Wilson_Harris
Wilson Pickett	http://en.wikipedia.org/wiki/Wilson_Pickett
Wilt Chamberlain	http://en.wikipedia.org/wiki/Wilt_Chamberlain
Wilton Persons	http://en.wikipedia.org/wiki/Wilton_Persons
Wim Wenders	http://en.wikipedia.org/wiki/Wim_Wenders
Winfield Scott	http://en.wikipedia.org/wiki/Winfield_Scott
Winfield Scott Hancock	http://en.wikipedia.org/wiki/Winfield_Scott_Hancock
Wings Hauser	http://en.wikipedia.org/wiki/Wings_Hauser
Wink Martindale	http://en.wikipedia.org/wiki/Wink_Martindale
Winnie Mandela	http://en.wikipedia.org/wiki/Winnie_Mandela
Winona Ryder	http://en.wikipedia.org/wiki/Winona_Ryder
Winslow Homer	http://en.wikipedia.org/wiki/Winslow_Homer
Winston Churchill	http://en.wikipedia.org/wiki/Winston_Churchill
Winston Churchill	http://en.wikipedia.org/wiki/Winston_Churchill_(novelist)
Winthrop Rockefeller	http://en.wikipedia.org/wiki/Winthrop_Rockefeller
Winthrop Sargent	http://en.wikipedia.org/wiki/Winthrop_Sargent
Wislawa Szymborska	http://en.wikipedia.org/wiki/Wislawa_Szymborska
Witold Lutoslawski	http://en.wikipedia.org/wiki/Witold_Lutoslawski
Wladyslaw Gomulka	http://en.wikipedia.org/wiki/Wladyslaw_Gomulka
Wojciech Jaruzelski	http://en.wikipedia.org/wiki/Wojciech_Jaruzelski
Wole Soyinka	http://en.wikipedia.org/wiki/Wole_Soyinka
Wolf Blitzer	http://en.wikipedia.org/wiki/Wolf_Blitzer
Wolfgang Amadeus Mozart	http://en.wikipedia.org/wiki/Wolfgang_Amadeus_Mozart
Wolfgang Amadeus Mozart	http://en.wikipedia.org/wiki/Wolfgang_Amadeus_Mozart
Wolfgang Capito	http://en.wikipedia.org/wiki/Wolfgang_Capito
Wolfgang Dauner	http://en.wikipedia.org/wiki/Wolfgang_Dauner
Wolfgang Ketterle	http://en.wikipedia.org/wiki/Wolfgang_Ketterle
Wolfgang Paul	http://en.wikipedia.org/wiki/Wolfgang_Paul
Wolfgang Pauli	http://en.wikipedia.org/wiki/Wolfgang_Pauli
Wolfgang Petersen	http://en.wikipedia.org/wiki/Wolfgang_Petersen
Wolfgang Preiss	http://en.wikipedia.org/wiki/Wolfgang_Preiss
Wolfgang Puck	http://en.wikipedia.org/wiki/Wolfgang_Puck
Wolfgang Reitherman	http://en.wikipedia.org/wiki/Wolfgang_Reitherman
Wolfgang Sch�uble	http://en.wikipedia.org/wiki/Wolfgang_Sch%E4uble
Wolfgang Sch�ssel	http://en.wikipedia.org/wiki/Wolfgang_Sch%FCssel
Wolfgang Sch�ssel	http://en.wikipedia.org/wiki/Wolfgang_Sch%FCssel
Wolfman Jack	http://en.wikipedia.org/wiki/Wolfman_Jack
Wolfram von Eschenbach	http://en.wikipedia.org/wiki/Wolfram_von_Eschenbach
Wonsuk Chin	http://en.wikipedia.org/wiki/Wonsuk_Chin
Wood Harris	http://en.wikipedia.org/wiki/Wood_Harris
Woodrow Wilson	http://en.wikipedia.org/wiki/Woodrow_Wilson
Woody Allen	http://en.wikipedia.org/wiki/Woody_Allen
Woody Guthrie	http://en.wikipedia.org/wiki/Woody_Guthrie
Woody Harrelson	http://en.wikipedia.org/wiki/Woody_Harrelson
Woody Herman	http://en.wikipedia.org/wiki/Woody_Herman
Woody Strode	http://en.wikipedia.org/wiki/Woody_Strode
Woody Woodmansey	http://en.wikipedia.org/wiki/Woody_Woodmansey
Wright Morris	http://en.wikipedia.org/wiki/Wright_Morris
Wrong Way Corrigan	http://en.wikipedia.org/wiki/Wrong_Way_Corrigan
Wu Yi	http://en.wikipedia.org/wiki/Wu_Yi
Wyatt Earp	http://en.wikipedia.org/wiki/Wyatt_Earp
Wyche Fowler, Jr.	http://en.wikipedia.org/wiki/Wyche_Fowler%2C_Jr.
Wyclef Jean	http://en.wikipedia.org/wiki/Wyclef_Jean
Wyndham Lewis	http://en.wikipedia.org/wiki/Wyndham_Lewis
Wynonna Judd	http://en.wikipedia.org/wiki/Wynonna_Judd
Wynton Marsalis	http://en.wikipedia.org/wiki/Wynton_Marsalis
X. J. Kennedy	http://en.wikipedia.org/wiki/X._J._Kennedy
Xanana Gusm�o	http://en.wikipedia.org/wiki/Xanana_Gusm%E3o
Xander Berkeley	http://en.wikipedia.org/wiki/Xander_Berkeley
Xavier Becerra	http://en.wikipedia.org/wiki/Xavier_Becerra
Xavier Cugat	http://en.wikipedia.org/wiki/Xavier_Cugat
Xaviera Hollander	http://en.wikipedia.org/wiki/Xaviera_Hollander
Xeni Jardin	http://en.wikipedia.org/wiki/Xeni_Jardin
Xerxes the Great	http://en.wikipedia.org/wiki/Xerxes_the_Great
Y. A. Tittle	http://en.wikipedia.org/wiki/Y._A._Tittle
Yahoo Serious	http://en.wikipedia.org/wiki/Yahoo_Serious
Yahya Jammeh	http://en.wikipedia.org/wiki/Yahya_Jammeh
Yakov Smirnoff	http://en.wikipedia.org/wiki/Yakov_Smirnoff
Yakubu Gowon	http://en.wikipedia.org/wiki/Yakubu_Gowon
Yamil Adorno	http://en.wikipedia.org/wiki/Yamil_Adorno
Yamila Diaz	http://en.wikipedia.org/wiki/Yamila_Diaz
Yancy Butler	http://en.wikipedia.org/wiki/Yancy_Butler
Yang Liwei	http://en.wikipedia.org/wiki/Yang_Liwei
Yang Shangkun	http://en.wikipedia.org/wiki/Yang_Shangkun
Yang Zhiya	http://en.wikipedia.org/wiki/Yang_Zhiya
Yaphet Kotto	http://en.wikipedia.org/wiki/Yaphet_Kotto
Yasmeen Ghauri	http://en.wikipedia.org/wiki/Yasmeen_Ghauri
Yasmin Le Bon	http://en.wikipedia.org/wiki/Yasmin_Le_Bon
Yasmin Qureshi	http://en.wikipedia.org/wiki/Yasmin_Qureshi
Yasmine Bleeth	http://en.wikipedia.org/wiki/Yasmine_Bleeth
Yasser Arafat	http://en.wikipedia.org/wiki/Yasser_Arafat
Yasuhiro Nakasone	http://en.wikipedia.org/wiki/Yasuhiro_Nakasone
Yasuzo Masumura	http://en.wikipedia.org/wiki/Yasuzo_Masumura
Yayi Boni	http://en.wikipedia.org/wiki/Yayi_Boni
Yeardley Smith	http://en.wikipedia.org/wiki/Yeardley_Smith
Yegor Ligachev	http://en.wikipedia.org/wiki/Yegor_Ligachev
Yehudi Menuhin	http://en.wikipedia.org/wiki/Yehudi_Menuhin
Yelena Bonner	http://en.wikipedia.org/wiki/Yelena_Bonner
Yelena Koreneva	http://en.wikipedia.org/wiki/Yelena_Koreneva
Yevgeny Primakov	http://en.wikipedia.org/wiki/Yevgeny_Primakov
Yevgeny Yevtushenko	http://en.wikipedia.org/wiki/Yevgeny_Yevtushenko
Yitzhak Rabin	http://en.wikipedia.org/wiki/Yitzhak_Rabin
Yitzhak Shamir	http://en.wikipedia.org/wiki/Yitzhak_Shamir
Yma Sumac	http://en.wikipedia.org/wiki/Yma_Sumac
Yngwie Malmsteen	http://en.wikipedia.org/wiki/Yngwie_Malmsteen
Yogi Berra	http://en.wikipedia.org/wiki/Yogi_Berra
Yoko Ono	http://en.wikipedia.org/wiki/Yoko_Ono
Yolanda Adams	http://en.wikipedia.org/wiki/Yolanda_Adams
Yordan Radichkov	http://en.wikipedia.org/wiki/Yordan_Radichkov
Yoshiro Mori	http://en.wikipedia.org/wiki/Yoshiro_Mori
Yotaro Kobayashi	http://en.wikipedia.org/wiki/Yotaro_Kobayashi
Young Buck	http://en.wikipedia.org/wiki/Young_Buck
Young Jeezy	http://en.wikipedia.org/wiki/Young_Jeezy
Young Jessie	http://en.wikipedia.org/wiki/Young_Jessie
Young MC	http://en.wikipedia.org/wiki/Young_MC
Young Vivian	http://en.wikipedia.org/wiki/Young_Vivian
Younghill Kang	http://en.wikipedia.org/wiki/Younghill_Kang
Yousaf Raza Gillani	http://en.wikipedia.org/wiki/Yousaf_Raza_Gillani
Yousuf Karsh	http://en.wikipedia.org/wiki/Yousuf_Karsh
Yoweri Museveni	http://en.wikipedia.org/wiki/Yoweri_Museveni
Yo-Yo Ma	http://en.wikipedia.org/wiki/Yo-Yo_Ma
Yuan T. Lee	http://en.wikipedia.org/wiki/Yuan_T._Lee
Yukihiro Matsumoto	http://en.wikipedia.org/wiki/Yukihiro_Matsumoto
Yukio Mishima	http://en.wikipedia.org/wiki/Yukio_Mishima
Yul Brynner	http://en.wikipedia.org/wiki/Yul_Brynner
Yuri Amano	http://en.wikipedia.org/wiki/Yuri_Amano
Yuri Andropov	http://en.wikipedia.org/wiki/Yuri_Andropov
Yuri Gagarin	http://en.wikipedia.org/wiki/Yuri_Gagarin
Yury Morozov	http://en.wikipedia.org/wiki/Yury_Morozov
Yusef Komunyakaa	http://en.wikipedia.org/wiki/Yusef_Komunyakaa
Yutake Ishinabe	http://en.wikipedia.org/wiki/Yutake_Ishinabe
Yuvraj Singh	http://en.wikipedia.org/wiki/Yuvraj_Singh
Yves Leterme	http://en.wikipedia.org/wiki/Yves_Leterme
Yves Montand	http://en.wikipedia.org/wiki/Yves_Montand
Yves Saint Laurent	http://en.wikipedia.org/wiki/Yves_Saint_Laurent_(designer)
Yvette Cooper	http://en.wikipedia.org/wiki/Yvette_Cooper
Yvette D. Clarke	http://en.wikipedia.org/wiki/Yvette_D._Clarke
Yvette Mimieux	http://en.wikipedia.org/wiki/Yvette_Mimieux
Yvonne Craig	http://en.wikipedia.org/wiki/Yvonne_Craig
Yvonne De Carlo	http://en.wikipedia.org/wiki/Yvonne_De_Carlo
Yvonne Dionne	http://en.wikipedia.org/wiki/Yvonne_Dionne
Yvonne Fovargue	http://en.wikipedia.org/wiki/Yvonne_Fovargue
Yvor Winters	http://en.wikipedia.org/wiki/Yvor_Winters
Zac Efron	http://en.wikipedia.org/wiki/Zac_Efron
Zac Goldsmith	http://en.wikipedia.org/wiki/Zac_Goldsmith
Zac Hanson	http://en.wikipedia.org/wiki/Zac_Hanson
Zacarias Moussaoui	http://en.wikipedia.org/wiki/Zacarias_Moussaoui
Zach Braff	http://en.wikipedia.org/wiki/Zach_Braff
Zach Galligan	http://en.wikipedia.org/wiki/Zach_Galligan
Zach Wamp	http://en.wikipedia.org/wiki/Zach_Wamp
Zachary Scott	http://en.wikipedia.org/wiki/Zachary_Scott
Zachary Taylor	http://en.wikipedia.org/wiki/Zachary_Taylor
Zachery Ty Bryan	http://en.wikipedia.org/wiki/Zachery_Ty_Bryan
Zack de la Rocha	http://en.wikipedia.org/wiki/Zack_de_la_Rocha
Zack Space	http://en.wikipedia.org/wiki/Zack_Space
Zakir Hussain	http://en.wikipedia.org/wiki/Zakir_Hussain_(musician)
Zakir Hussain	http://en.wikipedia.org/wiki/Zakir_Hussain_(politician)
Zakk Wylde	http://en.wikipedia.org/wiki/Zakk_Wylde
Zander Schloss	http://en.wikipedia.org/wiki/Zander_Schloss
Zane Grey	http://en.wikipedia.org/wiki/Zane_Grey
Zazu Pitts	http://en.wikipedia.org/wiki/Zazu_Pitts
Zbigniew Brzezinski	http://en.wikipedia.org/wiki/Zbigniew_Brzezinski
Zdzislaw Beksinski	http://en.wikipedia.org/wiki/Zdzislaw_Beksinski
Zebulon Pike	http://en.wikipedia.org/wiki/Zebulon_Pike
Zebulon Vance	http://en.wikipedia.org/wiki/Zebulon_Vance
Zeena Parkins	http://en.wikipedia.org/wiki/Zeena_Parkins
Zeenat Aman	http://en.wikipedia.org/wiki/Zeenat_Aman
Zeferino dos Prazeres	http://en.wikipedia.org/wiki/Zeferino_dos_Prazeres
Zelda Rubinstein	http://en.wikipedia.org/wiki/Zelda_Rubinstein
Zelimkhan Yandarbiyev	http://en.wikipedia.org/wiki/Zelimkhan_Yandarbiyev
Zell Miller	http://en.wikipedia.org/wiki/Zell_Miller
Zentani Muhammad az-Zentani	http://en.wikipedia.org/wiki/Zentani_Muhammad_az-Zentani
Zeppo Marx	http://en.wikipedia.org/wiki/Zeppo_Marx
Zero Mostel	http://en.wikipedia.org/wiki/Zero_Mostel
Zev Yaroslavsky	http://en.wikipedia.org/wiki/Zev_Yaroslavsky
Zhao Ziyang	http://en.wikipedia.org/wiki/Zhao_Ziyang
Zhelyu Zhelev	http://en.wikipedia.org/wiki/Zhelyu_Zhelev
Zhores I. Alferov	http://en.wikipedia.org/wiki/Zhores_I._Alferov
Zhou Enlai	http://en.wikipedia.org/wiki/Zhou_Enlai
Ziaur Rahman	http://en.wikipedia.org/wiki/Ziaur_Rahman
Ziggy Marley	http://en.wikipedia.org/wiki/Ziggy_Marley
Zigmantas Balcytis	http://en.wikipedia.org/wiki/Zigmantas_Balcytis
Zillur Rahman	http://en.wikipedia.org/wiki/Zillur_Rahman
Zine El Abidine Ben Ali	http://en.wikipedia.org/wiki/Zine_El_Abidine_Ben_Ali
Zin�dine Zidane	http://en.wikipedia.org/wiki/Zin%E9dine_Zidane
Ziyi Zhang	http://en.wikipedia.org/wiki/Ziyi_Zhang
Zo� Baird	http://en.wikipedia.org/wiki/Zo%EB_Baird
Zoe Caldwell	http://en.wikipedia.org/wiki/Zoe_Caldwell
Zoe Lofgren	http://en.wikipedia.org/wiki/Zoe_Lofgren
Zoe Zaldana	http://en.wikipedia.org/wiki/Zoe_Zaldana
Zolt�n Kod�ly	http://en.wikipedia.org/wiki/Zolt%E1n_Kod%E1ly
Zona Gale	http://en.wikipedia.org/wiki/Zona_Gale
Zooey Deschanel	http://en.wikipedia.org/wiki/Zooey_Deschanel
Zoogz Rift	http://en.wikipedia.org/wiki/Zoogz_Rift
Zora Neale Hurston	http://en.wikipedia.org/wiki/Zora_Neale_Hurston
Zoran Amar	http://en.wikipedia.org/wiki/Zoran_Amar
Zsa Zsa Gabor	http://en.wikipedia.org/wiki/Zsa_Zsa_Gabor
Zulfikar Ali Bhutto	http://en.wikipedia.org/wiki/Zulfikar_Ali_Bhutto
Zurab Nogaideli	http://en.wikipedia.org/wiki/Zurab_Nogaideli
Zviad Gamsakhurdia	http://en.wikipedia.org/wiki/Zviad_Gamsakhurdia
