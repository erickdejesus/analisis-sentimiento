Mike Marshall	Programing Genius
Jeff Catlin	Evil Slavedriver :)
