100% Natural
3d Lashes
5D Movie
Abito
Acapella
Accesorios Celulares
Accycel
Actinver
Acuario Mr. Tortus
Adidas
Adidas Originals
Adixxion Maak
Adolfo Dominguez
Adrenalina
Adventure
Aerom�xico
A�ropostale
Aerosoles
AG
Albaricoque Couture
Albertos
Alboa
Aldo
Aldo Conti
Aldo Conti Jr
Alfilo
All Sport
American Eagle
American Health
Amk
Anabel
Anel et Chuy
Anelli Joyas
ANELLO
Antigua
Antojitos Emy
Applebees
Aqua Terra
Arabiga
Arantza
Argentina  Express
Arnoldi
Arrachera House
Arte Egipcio
Artesan�as de Tabasco
Asadero Beef
A-Takear
Audio Mundo
Autolasa
Aviso Oportuno
AXA Seguros
Ay G�ey
Aysha
Azul Pastel
B fashion
Baby Creysi
Baby Panda
Baby Up
Baby Upscale
Bah�a Sport Gym
Bai Hao
Bamboo
Banamex
Banana Republic
Bancomer
Bancomer cajeros
Banorte
Bari
Barrio Tinto
Be Cool
Beauty Salon Marisol
Bebe
Beefer�s
Bejjani
Bell�sima
Benedetti�s Pizza
Bernardi Caffe
Bershka
Bestday
Betty�s Burgers
Bewasp
Bia Brazil
Big Bola
Bimba y Lola
Biopiel
Bistrot Sainz
Bizzarro
Blitzer accesorios
Blitzer Jeans
Blossom Spa
Blsk
Blu Lagoon
Bo & Co
Boba Shot
Bobois
Boga
Bogart
Bol Perinorte
Bonga Gym
Boston�s
Botanicus
Brantano
Bras y mucho m�s
BRUNO CORZA
Buchakas
Build-A-Bear Workshop
Bull Rider
Bunaday
Bunraku
Burger King
Burritos El Punto
Burritos Factory
Burro-T
C&A
Cablecom
Cablemas
Cablevisi�n
Cabo Grill
Caf� Central
Cafe Finca Santa Veracruz
Cafe Frappisimo
Caf� Jekemir
Caf� Mozart
Caf� Punta del Cielo
Caf� Society
California Pizza Kitchen
California Prime Rib
Calle Tijera
Calvin Klein
Calzedonia Intimissimi
Campanita
Camper
Candy
Candy Bar
Capa de Ozono
Capa de Ozono 2
Caramela
Carl�s Jr
Carlo Giovanni
Carlo Rossetti
Carnevali
Carnitas Esteban
Carnitas La Esperanza
Carranza y Carranza
Carter's
Casa Arles
Casa de las Lomas
Casa Ortiz
Casino Joker
Casino Life
Cassava Roots
CAT Telcel
Catalina Vargas
Celular Express
Cencel
Cencel 2
Centro de Atenci�n a Clientes Telcel
Centro de Belleza Maru Sol�s
Ceviche�s
Charly
Charro
Chicco
Chicken House & Salads
Chico�s
Chili�s
Chilim Balam
Chilo Flautas
China Express
China Inn
China Town
Chi-Palace
Christine
Chrysler
Chuy�s Barber Shop
CI Banco
Cielito Querido Caf�
Cinemex
Cin�polis
Citizen
Click Joyas
Cloe
Club Premier Aeromexico
Cocinas integrales HA
Cocinas Quetzal
Cocodrilo Green
Coiffure Sebastian
Colorspot
Coloso
Columbia
Comatemi
Comic
Comic Baby
Comicx
Comunicaci�n Royal
Confetty
Confite
Contempo
Continental Gallery
Converse
Cool
Cool Fashion
Coqueta y Audaz
Correa Zapater�as
Cortefiel
Costa Line
Costushop
Crabtree & Evelyn
Crepe Corner
Crepes & Waffles
Cristal Joyas
Crochet
Crocs
Cuadra
Cuidado con el Perro
Dairy Queen
Daniel Espinosa
Danya Spa
Darinka
Daylight Salads
De Chile Mole y Pozole
Decor�
Deli Crepas
Delizie
Demi Jeans
Dentalia
Deperlas
Depila-t
Destination Maternity
Devlyn
Devlyn Solare
Devotchka
Di Bari Pizzeria
Di� Essenza
Diamantes y Perlas
Dic&Co
Dicass Sports
Dico
Didactijuegos
Digital Zone
Dione
Distroller Butik
Diversiones Galex
Divertido
Dk Boutique
Do&Be
Dockers
Dolce Mondo
Domino�s Pizza
Donal Top Salon
Dormimundo
Dorothy Gara
Dorothy Gaynor
Dorothy Gaynor 2
DP Street
Dportenis
dpstreet
Dry Clean USA
Dulcer�a Chile Nitz�
Dulcer�a D'Leal
D-U�as
DUO
Dynasty Chinese Food
Eclipse
Eclipse Plus
Ecobike
El Atico
El Corte Ingl�s
El Fog�n
El Galp�n Argentino
El Garabato
El Globo
El Jaripeo
El Mexicano
El ote
El P�ndulo
El Port�n
El Tinacal
El Torito
El Viajero del Norte
Elegance
Elite Lockers
Ellie Boutique
Elote Real
Emotion Casino
Emwa
Emyco
Enrique Bricker
Ensaladetti
Epicland
Erez
Ermenegildo Zegna
Es Coiffeurs
Escrupulos
Estaci�n del tren
Estefan�a Duarte Plata
Est�tica Bogus
Etam
Eternity Diamonds
Europiel Laser Center
Evoll�ser
Exotic
Exotica
Expo Plaza
Expressiones
Fabricas de Francia
Fabrizio
Faces
Fans Shop
Farmacia Benavides
Farmacias Yza
Fashionalia
Ferriano
Ferrioni
Ferrioni N1
Festivities Yayis
Fg Gaud�
Fiore Gelato
Fiorentina
Fitness Station
Flamin Wings
Flavio Gatto
Flexi
Florsheim
Fonda Santa Clara
Fonix distribuidor autorizado Telcel
Forever 21
Forever Teens
Foto F�cil
Fracmar
Franco Cuadra
Fresa
Friso
Frutiyogurth
Fullsand
Fundaci�n Dond�
Furor
G Candila
G.I in Style
Galer�as Florencia
Galer�as Rojas
Game Planet
Gandhi
Gap
Garabatos
Gelateria Italiana
Gelato
Georgie Boy
Georgie Boy 2
Giannino' s
Gigi�s Pizzeria
Giolini
Giovanni�s
Girls
Glazier
Gloria Jeans
GNC
Go Beauty
Goc
Gonher
Gonia
Gorditas Do�a Tota
Green Grass
Gre�itas
Guayaberass
Guess
Gula
Gushto
Guvier
H&M
H�agen Dazs
Hang Ten
Hawaiian Paradise
Heaven
Heaven PB
Helados Dairy Queen
Helados Nutrisa
Helados Santa Clara
Helados Sultana
Heroes Restaurant & Bar
Hey Fitness
Hidalgo
High Life
High Street
Hill�s
Holanda
Hotel Fiesta Inn
HP
HP store
HSBC
Hugo Boss
Hurley
Huun Libros & Lounge
Ice Gallerie
ICEDOME
Ichiban
If
Illro
Imaginarium
In Moda
Inbursa
Ingenia Muebles
Innova Sport
Innvictus
Insalades
Insoportablemente Argentino
Intempo
Interlingua
Isadora
Ishop
It
Italia Joyas
Italian Coffee
Italian Steak House
Italianni�s
Italiato
Italimo
Iusacell
Ivonne
Ivory Tours
Ixe Banco
Jarking
Jean Pierre
Jeans Beronna
Jeff de Bruges
Jobama
Johnny Rockets
Johnston & Murphy
Jollpat
Joyer�a Ruiz Hermanos
Joyer�as Luna
Juguetibici
Juguetron
Julio
Julio Cepeda
Julio Rocha
Juniors Coiffure
Just Kids
Karol�s Gift Shop
Karukay
Kauffman
Kensao
Keten
Key Di Ci
KFC
Kids Star
Kiehl's
Kiko Donas
Kingbird
Kipling
Knova
Koaj
Kokopao
Komacy
K-rime Collection
Krispy Kreme
Kukis by Maru
Kurian
Kush
L�Occitane
La Baguette
La Blanquita
La bonita
La Caba�a
La Callana
La Canasta
La Casa de los Rompecabezas
La casa del buen marisco
La Casa del Fumador
La Casa del Pastor
La Ciudad de Colima
La Crepa
La Creper�a
La Cupcakeria
La Esmeralda
La Europea
La Fe
La Fundidora
La Milagresa
La Norte�a
La Oriental
La Poupe�
La Ranita
La Spezia
Lacoste
Lacoste accesorios
Las Alitas
Las Juanas Torter�a
Lavander�a Ahucast
Lavoro
Le Boom To
Le Sport Sac
Lefties
Levi�s
Lia Bose
Libreria Dante
Librer�a de la Mancha
Librer�a La Ventana
Lieb Tobacco
Lila
Lilia Godinez
Lily Pot
Linda Only Nails
Lineas
Little Closet
Liverpool
Liverpool Motos
Liverpool Restaurante
Liz Minelli
Llantas Royal
Lob
Lob Footwear
Lobby
Lobo Solo
Lombok Exotic Touch
London Styles
Long Cheng
Loops & Coffee
Los Bisquets Bisquets Obreg�n
Los de Pescado
Los Trompos
Lux Sport
Mabel
Mac
Mac Store
Magic Trek
Maison Kayser
Malib�
Mama M�a
Mando�s
Mango
Marco Viali
Maria Isabel
MARIKARLI
Mario Hernandez
Marsel
Mart�
M�s Visi�n
Mascotas Leo�s
Maskota
Massimo Dutti
Max Mara
Mc Donald�s
McDonald�s
MCO
Mea Culpa
Melendez Grill
Men�s Factory
Men�s Fashion
Merrell
Miberth
Michel Domit
Michelle
Mineralia
Mistertennis
Mixup
Miyako
Mobo
Mobo Shop
Moderna Sport
Moditelas
Monas y Monitos
Mont Blanc
Montecassino
Moon Jeans
Mora Azul
Morrikos
Motosport
Movistar
Moyo
Mr. Sushi
Muebles Dico
Mujer Bonita
Mundo Feliz
Mundo Helado
Mundo Odontol�gico
Mundo Peque
Musas
Muzza
Muzza Zapater�a
Mystic
Nana Pancha
Narda
Nathan�s
Natural
Natural Scents
Naturale�s
Naturhouse
Nespresso
Nestle
Neve Gelato
New Gym
Nextel
Nicholas
Nike
Nike Store
N�na Ferr�
Nine West
Novart Boutique
Nuny's Yogurt
Nutrisa
Oh lala
Oh! Interiorismo Contempor�neo
Okey
Omnia Boutique
Onix
Only Nail
Opp�s Jeans
Optica Americana
Optica Mirely
Opticas Am�rica
Opticas Lux
Optikal & Krono Shop
Oriental Wok
Orios Boutique
Oro y Plata de Colecci�n
Orthodontics Center of America
Oshkosh
Oxido
Oxxo
Oysho
P.F. Chang�s China Bistro
P.S. by A�ropostale
Palacio de Hierro
Palacio de Hierro - Restaurante
Pampa y Tango
Pandora
Pao Lee
Papillon
Papo�s Shoes
Parfums Rachelle
Parrilla del Charro
Paseli
Passion
Pasteler�a Americana
Pasteler�a Lolita
Patrice
Patrotur
Paul & Shark
Pavi Italy
Paws
Penguin
People in Red
Pepe Jeans
Pepper�s
Perfect Choice
Perugia
Petland
PG Beauty
Phiten
Phone City
Photofolio
Pia Makart
Piacenza Ristorante
Piccolo Mondo
Pick a Sandwich
Piedi Carino
Piel de Plata
Pikolinos
Piky Accessories
Pirma
Pizza Amore
Pizza Hut
Pizza Hut Restaurante
Pizzer�a Di Bari
Pizzer�a Romana
Pizzeria y tacos de mariscos Marea
Pizzeta
Plata de Taxco
Platax & Co
Play Circus
Play City
Play Time
Playland
PODO CARE
Polo Club
Polo Sur
Ponte Almeja
Pop Atelier
Pop Bar
Prada
Presta Prenda  Banco Azteca
Professional Cycling
Prostyle
Pull and Bear
Puma
Puma Time
Punto Muerto
Puro Pollo
Qing Dao
Quarry
Queen
Quick Cut
Quiksilver
Quilmes
Quinto Piso
Quiznos
Quiznos Restaurante
R Julian
R. Picard
Radio Shack
Rafa Velasco Estilista
Ram
Rana�s
Recorcholis
Red Mango
Regalos El Chapul�n
Rin Rin Pizza
Rinc�n Chino
Rio Grande
River's System
Robert�s
Rock Hampton
Rossati
Rous the Shoe Boutique
Royal Prestige
Rudos
Run Freaks
Sahari�s
Sally Beauty Supply
Salomon
Samsonite
San Cerdito
Sanborns
Sandra
Sanrio Smiles
Sanrio Surprises
Santa Clara
Santander Serf�n
Santangel
Sayori
Sbarro
Scappino
Scappino 2
Schiaparelli
Scotiabank Inverlat
Sears
Sebastian
Sebastian Lashes
Segafredo
Servitime
Sexy Jeans
Sfera
Shari Maki
Shasa
SHASTRA
Shi Wei Xian
Shoe Xotica
Silvia Carnevali
Sirloin Stockade
Sisters Forever
Sixties
Skechers
Skin Care Kopay
Slim Center
Slinky
Small Animals
Smart Fit
Smartfone
Snack
Snob Bistro
Solaris
Sole
Soley
Sony Store
Soriana
Sorpelle
Sorrento
Spa Sebasti�n
Spalding
Specialized
Sportia
Sportif
Sportortas
Springfield
Squalo
St Even
Starbucks
Stellari
Stephanie Ascencio
Steren
Steren Shop
Sterling
Steve Madden
Stilisimo
Stop
Storm Extreme
Storm Gotcha
Stradivarius
Stuarts
Studio
Studio F
Studio Hair Saloon
Stylo
Subway
Subway Restaurante
Sunglass Hut
S�per Salads
Surman
Sushi Itto
Sushi Roll
Sushi Roll Restaurante
Sushi Salads
Swarovski
Swatch
Taco Beef
Taco Inn
Taco Maran
TAF
Tamaris
Tane
Tapioca House
Taquitos de Pm
Tara Brooch
Tarocco
Tea & Coffee House
Ted Kenton
Teddy Mountain
Telcel
Tempo
Tennis Star
Teriyaki San
Texas Ribs
Thai & Japan
The Best House
The Body Shop
The Boss Place
The Coffee Time
The Italian Coffee
The Met
The Nail Corner
The Urban Corner
Thrifty
Tierra del fuego
Tio Taco
Todo Moda
Todo para sus pies
Toks
Tommy Hilfiger
Topp's
Tops & Bottoms
Tortas.com
Torton�s
Toscano
Totto
Tous
Toxic
Trender
Trenes Insurgentes
Trini
trueKDS
TT Blues
Tucan�
Tufan Tapetes
Turin
TV Tiendas
Two Par Kids
U Adolfo Dominguez
Unagui
United Airlines
United Colors Of Benetton
U�as Finas
U�as Norma
Ups Regalos
UPS!
Urban Looks
Utopia
Valentina
Vallarta Fitness
Vanita
Vanity
Vans
Vaso Loko
Veerkamp
Veika
Vela piel
Velatti Muebles
Vell�simo
Vertiche
Very Sexy
Veterinaria Mascotas Koala
V�a Rep�blica
Via Uno
Viajes Intermex
Viajes Palacio
Viajes Tabasco
Vicky Form
Victoria Piel y Mas
Victoria�s Secret
Vida Marina
Vilebrequin
Violeta by Mango
VIP Global Solutions
Vip�s
Vira Vira
Visi�n �ptica
Visual Tendence
Vittorio Forti
Vohua
Walking Toes
Wall�s BabersShop
Walmart
wb
Wendy�s
Wings Army
Women� Secret
Woods
Xerox
Xunxes
Yak Sports & Books
Yanina
Yaska
Yeno�
Yogen fruz
Yokiro Sushi
Yomi Wok
Yomood
Yong Chang
Yozen
Yumorama
Yves Rocher
Zara
Zara Home
Zara N1
Zingara
Zoe Collection
Zurich